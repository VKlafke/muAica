library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.muAica_pkg.all;

entity muAica_tb is
end entity muAica_tb;

architecture behavior of muAica_tb is

  -- processor top module component
  COMPONENT muAica is
    port (
      clk       : in    std_logic;
      rst_bt    : in    std_logic;
      port_io   : inout std_logic_vector (n-1 downto 0); -- configurable IO port
      tx        : out std_logic;
	    rx: in std_logic
    );
  end COMPONENT muAica;

  -- System clock and reset
  signal  clk   : std_logic;
  signal  rst_bt: std_logic;

  constant half_period : time := 10 ns; -- 50 MHZ

  signal  intr_sig : std_logic;
  signal  port_io_sig  : std_logic_vector (n-1 downto 0); -- interface with microcontroller port

  signal tx_s : std_logic; -- tx signal
  signal rx_s : std_logic;

  signal tx_dv : std_logic;
  signal tx_active_s : std_logic;
  signal tx_done :std_logic;
  signal data_tx : std_logic_vector(7 downto 0);

begin

  -- Clock process: 100 MHz
  signal_clk : process
  begin
    clk <= '0'; wait for half_period;
    loop
      clk <= '1'; wait for half_period;
      clk <= '0'; wait for half_period;
    end loop;
  end process signal_clk;

  -- Clock
  rst_button : process -- debounce should be disabled inside 'aica/bt_debounce' (stability time ~0)
  begin
    rst_bt <= '0'; wait for 100 ns;
    loop
      rst_bt <= '1'; wait for 50 ns;
      rst_bt <= '0'; wait for 20 sec;
      rst_bt <= '1'; wait for 100 ns;
      rst_bt <= '0'; wait for 10 sec;
    end loop;
  end process rst_button;

-- Port Map
  MICRO_AICA: muAica
  port map(
    clk     => clk,
    rst_bt  => rst_bt,
    port_io => port_io_sig,
    tx      => tx_s,
	  rx		=> rx_s
  );
  
 -- rx_s <= '0';

  -- Send data to rx
  TX_DATA_SEND: entity work.UART_TX_v1
  port map(
    i_Clk       => clk,
    i_TX_DV     => tx_dv,
    i_TX_Byte   => data_tx,
    o_TX_Active => tx_active_s,
    o_TX_Serial => rx_s,
    o_TX_Done   => tx_done
  );

-- VHDL for data_tx:
data_tx <= x"00" after 0 ns,
x"00" after 11000 ns,
x"09" after 22000 ns,
x"AC" after 33000 ns,
x"17" after 44000 ns,
x"21" after 55000 ns,
x"00" after 66000 ns,
x"00" after 77000 ns,
x"13" after 88000 ns,
x"01" after 99000 ns,
x"01" after 110000 ns,
x"43" after 121000 ns,
x"13" after 132000 ns,
x"01" after 143000 ns,
x"C1" after 154000 ns,
x"FF" after 165000 ns,
x"23" after 176000 ns,
x"20" after 187000 ns,
x"11" after 198000 ns,
x"00" after 209000 ns,
x"37" after 220000 ns,
x"1F" after 231000 ns,
x"00" after 242000 ns,
x"00" after 253000 ns,
x"13" after 264000 ns,
x"0F" after 275000 ns,
x"0F" after 286000 ns,
x"80" after 297000 ns,
x"73" after 308000 ns,
x"20" after 319000 ns,
x"4F" after 330000 ns,
x"30" after 341000 ns,
x"73" after 352000 ns,
x"60" after 363000 ns,
x"44" after 374000 ns,
x"30" after 385000 ns,
x"73" after 396000 ns,
x"60" after 407000 ns,
x"04" after 418000 ns,
x"30" after 429000 ns,
x"73" after 440000 ns,
x"10" after 451000 ns,
x"10" after 462000 ns,
x"34" after 473000 ns,
x"73" after 484000 ns,
x"10" after 495000 ns,
x"20" after 506000 ns,
x"34" after 517000 ns,
x"EF" after 528000 ns,
x"00" after 539000 ns,
x"50" after 550000 ns,
x"01" after 561000 ns,
x"83" after 572000 ns,
x"20" after 583000 ns,
x"01" after 594000 ns,
x"00" after 605000 ns,
x"13" after 616000 ns,
x"01" after 627000 ns,
x"41" after 638000 ns,
x"00" after 649000 ns,
x"67" after 660000 ns,
x"80" after 671000 ns,
x"00" after 682000 ns,
x"00" after 693000 ns,
x"93" after 704000 ns,
x"08" after 715000 ns,
x"10" after 726000 ns,
x"00" after 737000 ns,
x"73" after 748000 ns,
x"00" after 759000 ns,
x"00" after 770000 ns,
x"00" after 781000 ns,
x"67" after 792000 ns,
x"80" after 803000 ns,
x"00" after 814000 ns,
x"00" after 825000 ns,
x"93" after 836000 ns,
x"08" after 847000 ns,
x"30" after 858000 ns,
x"00" after 869000 ns,
x"73" after 880000 ns,
x"00" after 891000 ns,
x"00" after 902000 ns,
x"00" after 913000 ns,
x"67" after 924000 ns,
x"80" after 935000 ns,
x"00" after 946000 ns,
x"00" after 957000 ns,
x"93" after 968000 ns,
x"08" after 979000 ns,
x"40" after 990000 ns,
x"00" after 1001000 ns,
x"73" after 1012000 ns,
x"00" after 1023000 ns,
x"00" after 1034000 ns,
x"00" after 1045000 ns,
x"67" after 1056000 ns,
x"80" after 1067000 ns,
x"00" after 1078000 ns,
x"00" after 1089000 ns,
x"93" after 1100000 ns,
x"08" after 1111000 ns,
x"50" after 1122000 ns,
x"00" after 1133000 ns,
x"73" after 1144000 ns,
x"00" after 1155000 ns,
x"00" after 1166000 ns,
x"00" after 1177000 ns,
x"67" after 1188000 ns,
x"80" after 1199000 ns,
x"00" after 1210000 ns,
x"00" after 1221000 ns,
x"93" after 1232000 ns,
x"08" after 1243000 ns,
x"A0" after 1254000 ns,
x"00" after 1265000 ns,
x"73" after 1276000 ns,
x"00" after 1287000 ns,
x"00" after 1298000 ns,
x"00" after 1309000 ns,
x"67" after 1320000 ns,
x"80" after 1331000 ns,
x"00" after 1342000 ns,
x"00" after 1353000 ns,
x"93" after 1364000 ns,
x"08" after 1375000 ns,
x"B0" after 1386000 ns,
x"00" after 1397000 ns,
x"73" after 1408000 ns,
x"00" after 1419000 ns,
x"00" after 1430000 ns,
x"00" after 1441000 ns,
x"67" after 1452000 ns,
x"80" after 1463000 ns,
x"00" after 1474000 ns,
x"00" after 1485000 ns,
x"93" after 1496000 ns,
x"08" after 1507000 ns,
x"C0" after 1518000 ns,
x"00" after 1529000 ns,
x"73" after 1540000 ns,
x"00" after 1551000 ns,
x"00" after 1562000 ns,
x"00" after 1573000 ns,
x"67" after 1584000 ns,
x"80" after 1595000 ns,
x"00" after 1606000 ns,
x"00" after 1617000 ns,
x"93" after 1628000 ns,
x"08" after 1639000 ns,
x"D0" after 1650000 ns,
x"00" after 1661000 ns,
x"73" after 1672000 ns,
x"00" after 1683000 ns,
x"00" after 1694000 ns,
x"00" after 1705000 ns,
x"67" after 1716000 ns,
x"80" after 1727000 ns,
x"00" after 1738000 ns,
x"00" after 1749000 ns,
x"93" after 1760000 ns,
x"08" after 1771000 ns,
x"E0" after 1782000 ns,
x"00" after 1793000 ns,
x"73" after 1804000 ns,
x"00" after 1815000 ns,
x"00" after 1826000 ns,
x"00" after 1837000 ns,
x"67" after 1848000 ns,
x"80" after 1859000 ns,
x"00" after 1870000 ns,
x"00" after 1881000 ns,
x"93" after 1892000 ns,
x"08" after 1903000 ns,
x"F0" after 1914000 ns,
x"00" after 1925000 ns,
x"73" after 1936000 ns,
x"00" after 1947000 ns,
x"00" after 1958000 ns,
x"00" after 1969000 ns,
x"67" after 1980000 ns,
x"80" after 1991000 ns,
x"00" after 2002000 ns,
x"00" after 2013000 ns,
x"93" after 2024000 ns,
x"08" after 2035000 ns,
x"00" after 2046000 ns,
x"01" after 2057000 ns,
x"73" after 2068000 ns,
x"00" after 2079000 ns,
x"00" after 2090000 ns,
x"00" after 2101000 ns,
x"67" after 2112000 ns,
x"80" after 2123000 ns,
x"00" after 2134000 ns,
x"00" after 2145000 ns,
x"13" after 2156000 ns,
x"01" after 2167000 ns,
x"81" after 2178000 ns,
x"FE" after 2189000 ns,
x"23" after 2200000 ns,
x"2A" after 2211000 ns,
x"81" after 2222000 ns,
x"00" after 2233000 ns,
x"13" after 2244000 ns,
x"04" after 2255000 ns,
x"81" after 2266000 ns,
x"01" after 2277000 ns,
x"23" after 2288000 ns,
x"26" after 2299000 ns,
x"A4" after 2310000 ns,
x"FE" after 2321000 ns,
x"83" after 2332000 ns,
x"27" after 2343000 ns,
x"C4" after 2354000 ns,
x"FE" after 2365000 ns,
x"23" after 2376000 ns,
x"2A" after 2387000 ns,
x"F4" after 2398000 ns,
x"FE" after 2409000 ns,
x"6F" after 2420000 ns,
x"00" after 2431000 ns,
x"00" after 2442000 ns,
x"01" after 2453000 ns,
x"83" after 2464000 ns,
x"27" after 2475000 ns,
x"44" after 2486000 ns,
x"FF" after 2497000 ns,
x"93" after 2508000 ns,
x"87" after 2519000 ns,
x"17" after 2530000 ns,
x"00" after 2541000 ns,
x"23" after 2552000 ns,
x"2A" after 2563000 ns,
x"F4" after 2574000 ns,
x"FE" after 2585000 ns,
x"83" after 2596000 ns,
x"27" after 2607000 ns,
x"44" after 2618000 ns,
x"FF" after 2629000 ns,
x"83" after 2640000 ns,
x"C7" after 2651000 ns,
x"07" after 2662000 ns,
x"00" after 2673000 ns,
x"E3" after 2684000 ns,
x"96" after 2695000 ns,
x"07" after 2706000 ns,
x"FE" after 2717000 ns,
x"03" after 2728000 ns,
x"27" after 2739000 ns,
x"44" after 2750000 ns,
x"FF" after 2761000 ns,
x"83" after 2772000 ns,
x"27" after 2783000 ns,
x"C4" after 2794000 ns,
x"FE" after 2805000 ns,
x"B3" after 2816000 ns,
x"07" after 2827000 ns,
x"F7" after 2838000 ns,
x"40" after 2849000 ns,
x"13" after 2860000 ns,
x"85" after 2871000 ns,
x"07" after 2882000 ns,
x"00" after 2893000 ns,
x"03" after 2904000 ns,
x"24" after 2915000 ns,
x"41" after 2926000 ns,
x"01" after 2937000 ns,
x"13" after 2948000 ns,
x"01" after 2959000 ns,
x"81" after 2970000 ns,
x"01" after 2981000 ns,
x"67" after 2992000 ns,
x"80" after 3003000 ns,
x"00" after 3014000 ns,
x"00" after 3025000 ns,
x"13" after 3036000 ns,
x"01" after 3047000 ns,
x"81" after 3058000 ns,
x"FE" after 3069000 ns,
x"23" after 3080000 ns,
x"2A" after 3091000 ns,
x"81" after 3102000 ns,
x"00" after 3113000 ns,
x"13" after 3124000 ns,
x"04" after 3135000 ns,
x"81" after 3146000 ns,
x"01" after 3157000 ns,
x"23" after 3168000 ns,
x"26" after 3179000 ns,
x"A4" after 3190000 ns,
x"FE" after 3201000 ns,
x"23" after 3212000 ns,
x"24" after 3223000 ns,
x"B4" after 3234000 ns,
x"FE" after 3245000 ns,
x"23" after 3256000 ns,
x"2A" after 3267000 ns,
x"04" after 3278000 ns,
x"FE" after 3289000 ns,
x"6F" after 3300000 ns,
x"00" after 3311000 ns,
x"00" after 3322000 ns,
x"03" after 3333000 ns,
x"03" after 3344000 ns,
x"27" after 3355000 ns,
x"84" after 3366000 ns,
x"FE" after 3377000 ns,
x"93" after 3388000 ns,
x"07" after 3399000 ns,
x"17" after 3410000 ns,
x"00" after 3421000 ns,
x"23" after 3432000 ns,
x"24" after 3443000 ns,
x"F4" after 3454000 ns,
x"FE" after 3465000 ns,
x"83" after 3476000 ns,
x"27" after 3487000 ns,
x"C4" after 3498000 ns,
x"FE" after 3509000 ns,
x"93" after 3520000 ns,
x"86" after 3531000 ns,
x"17" after 3542000 ns,
x"00" after 3553000 ns,
x"23" after 3564000 ns,
x"26" after 3575000 ns,
x"D4" after 3586000 ns,
x"FE" after 3597000 ns,
x"03" after 3608000 ns,
x"47" after 3619000 ns,
x"07" after 3630000 ns,
x"00" after 3641000 ns,
x"23" after 3652000 ns,
x"80" after 3663000 ns,
x"E7" after 3674000 ns,
x"00" after 3685000 ns,
x"83" after 3696000 ns,
x"27" after 3707000 ns,
x"44" after 3718000 ns,
x"FF" after 3729000 ns,
x"93" after 3740000 ns,
x"87" after 3751000 ns,
x"17" after 3762000 ns,
x"00" after 3773000 ns,
x"23" after 3784000 ns,
x"2A" after 3795000 ns,
x"F4" after 3806000 ns,
x"FE" after 3817000 ns,
x"83" after 3828000 ns,
x"27" after 3839000 ns,
x"84" after 3850000 ns,
x"FE" after 3861000 ns,
x"83" after 3872000 ns,
x"C7" after 3883000 ns,
x"07" after 3894000 ns,
x"00" after 3905000 ns,
x"E3" after 3916000 ns,
x"96" after 3927000 ns,
x"07" after 3938000 ns,
x"FC" after 3949000 ns,
x"83" after 3960000 ns,
x"27" after 3971000 ns,
x"C4" after 3982000 ns,
x"FE" after 3993000 ns,
x"23" after 4004000 ns,
x"80" after 4015000 ns,
x"07" after 4026000 ns,
x"00" after 4037000 ns,
x"83" after 4048000 ns,
x"27" after 4059000 ns,
x"44" after 4070000 ns,
x"FF" after 4081000 ns,
x"13" after 4092000 ns,
x"85" after 4103000 ns,
x"07" after 4114000 ns,
x"00" after 4125000 ns,
x"03" after 4136000 ns,
x"24" after 4147000 ns,
x"41" after 4158000 ns,
x"01" after 4169000 ns,
x"13" after 4180000 ns,
x"01" after 4191000 ns,
x"81" after 4202000 ns,
x"01" after 4213000 ns,
x"67" after 4224000 ns,
x"80" after 4235000 ns,
x"00" after 4246000 ns,
x"00" after 4257000 ns,
x"13" after 4268000 ns,
x"01" after 4279000 ns,
x"81" after 4290000 ns,
x"FD" after 4301000 ns,
x"23" after 4312000 ns,
x"22" after 4323000 ns,
x"81" after 4334000 ns,
x"02" after 4345000 ns,
x"13" after 4356000 ns,
x"04" after 4367000 ns,
x"81" after 4378000 ns,
x"02" after 4389000 ns,
x"23" after 4400000 ns,
x"2E" after 4411000 ns,
x"A4" after 4422000 ns,
x"FC" after 4433000 ns,
x"23" after 4444000 ns,
x"2C" after 4455000 ns,
x"B4" after 4466000 ns,
x"FC" after 4477000 ns,
x"B7" after 4488000 ns,
x"17" after 4499000 ns,
x"00" after 4510000 ns,
x"00" after 4521000 ns,
x"93" after 4532000 ns,
x"87" after 4543000 ns,
x"87" after 4554000 ns,
x"85" after 4565000 ns,
x"83" after 4576000 ns,
x"A5" after 4587000 ns,
x"07" after 4598000 ns,
x"00" after 4609000 ns,
x"03" after 4620000 ns,
x"A6" after 4631000 ns,
x"47" after 4642000 ns,
x"00" after 4653000 ns,
x"83" after 4664000 ns,
x"A6" after 4675000 ns,
x"87" after 4686000 ns,
x"00" after 4697000 ns,
x"03" after 4708000 ns,
x"A7" after 4719000 ns,
x"C7" after 4730000 ns,
x"00" after 4741000 ns,
x"23" after 4752000 ns,
x"22" after 4763000 ns,
x"B4" after 4774000 ns,
x"FE" after 4785000 ns,
x"23" after 4796000 ns,
x"24" after 4807000 ns,
x"C4" after 4818000 ns,
x"FE" after 4829000 ns,
x"23" after 4840000 ns,
x"26" after 4851000 ns,
x"D4" after 4862000 ns,
x"FE" after 4873000 ns,
x"23" after 4884000 ns,
x"28" after 4895000 ns,
x"E4" after 4906000 ns,
x"FE" after 4917000 ns,
x"83" after 4928000 ns,
x"C7" after 4939000 ns,
x"07" after 4950000 ns,
x"01" after 4961000 ns,
x"23" after 4972000 ns,
x"0A" after 4983000 ns,
x"F4" after 4994000 ns,
x"FE" after 5005000 ns,
x"83" after 5016000 ns,
x"27" after 5027000 ns,
x"84" after 5038000 ns,
x"FD" after 5049000 ns,
x"93" after 5060000 ns,
x"D7" after 5071000 ns,
x"47" after 5082000 ns,
x"40" after 5093000 ns,
x"93" after 5104000 ns,
x"F7" after 5115000 ns,
x"F7" after 5126000 ns,
x"00" after 5137000 ns,
x"93" after 5148000 ns,
x"87" after 5159000 ns,
x"87" after 5170000 ns,
x"FF" after 5181000 ns,
x"B3" after 5192000 ns,
x"87" after 5203000 ns,
x"87" after 5214000 ns,
x"00" after 5225000 ns,
x"03" after 5236000 ns,
x"C7" after 5247000 ns,
x"C7" after 5258000 ns,
x"FE" after 5269000 ns,
x"83" after 5280000 ns,
x"27" after 5291000 ns,
x"C4" after 5302000 ns,
x"FD" after 5313000 ns,
x"23" after 5324000 ns,
x"80" after 5335000 ns,
x"E7" after 5346000 ns,
x"00" after 5357000 ns,
x"83" after 5368000 ns,
x"27" after 5379000 ns,
x"84" after 5390000 ns,
x"FD" after 5401000 ns,
x"13" after 5412000 ns,
x"F7" after 5423000 ns,
x"F7" after 5434000 ns,
x"00" after 5445000 ns,
x"83" after 5456000 ns,
x"27" after 5467000 ns,
x"C4" after 5478000 ns,
x"FD" after 5489000 ns,
x"93" after 5500000 ns,
x"87" after 5511000 ns,
x"17" after 5522000 ns,
x"00" after 5533000 ns,
x"13" after 5544000 ns,
x"07" after 5555000 ns,
x"87" after 5566000 ns,
x"FF" after 5577000 ns,
x"33" after 5588000 ns,
x"07" after 5599000 ns,
x"87" after 5610000 ns,
x"00" after 5621000 ns,
x"03" after 5632000 ns,
x"47" after 5643000 ns,
x"C7" after 5654000 ns,
x"FE" after 5665000 ns,
x"23" after 5676000 ns,
x"80" after 5687000 ns,
x"E7" after 5698000 ns,
x"00" after 5709000 ns,
x"83" after 5720000 ns,
x"27" after 5731000 ns,
x"C4" after 5742000 ns,
x"FD" after 5753000 ns,
x"93" after 5764000 ns,
x"87" after 5775000 ns,
x"27" after 5786000 ns,
x"00" after 5797000 ns,
x"23" after 5808000 ns,
x"80" after 5819000 ns,
x"07" after 5830000 ns,
x"00" after 5841000 ns,
x"93" after 5852000 ns,
x"07" after 5863000 ns,
x"20" after 5874000 ns,
x"00" after 5885000 ns,
x"13" after 5896000 ns,
x"85" after 5907000 ns,
x"07" after 5918000 ns,
x"00" after 5929000 ns,
x"03" after 5940000 ns,
x"24" after 5951000 ns,
x"41" after 5962000 ns,
x"02" after 5973000 ns,
x"13" after 5984000 ns,
x"01" after 5995000 ns,
x"81" after 6006000 ns,
x"02" after 6017000 ns,
x"67" after 6028000 ns,
x"80" after 6039000 ns,
x"00" after 6050000 ns,
x"00" after 6061000 ns,
x"13" after 6072000 ns,
x"01" after 6083000 ns,
x"01" after 6094000 ns,
x"FC" after 6105000 ns,
x"23" after 6116000 ns,
x"2E" after 6127000 ns,
x"81" after 6138000 ns,
x"02" after 6149000 ns,
x"13" after 6160000 ns,
x"04" after 6171000 ns,
x"01" after 6182000 ns,
x"04" after 6193000 ns,
x"23" after 6204000 ns,
x"22" after 6215000 ns,
x"A4" after 6226000 ns,
x"FC" after 6237000 ns,
x"23" after 6248000 ns,
x"20" after 6259000 ns,
x"B4" after 6270000 ns,
x"FC" after 6281000 ns,
x"23" after 6292000 ns,
x"2A" after 6303000 ns,
x"04" after 6314000 ns,
x"FE" after 6325000 ns,
x"23" after 6336000 ns,
x"26" after 6347000 ns,
x"04" after 6358000 ns,
x"FE" after 6369000 ns,
x"83" after 6380000 ns,
x"27" after 6391000 ns,
x"04" after 6402000 ns,
x"FC" after 6413000 ns,
x"93" after 6424000 ns,
x"D7" after 6435000 ns,
x"F7" after 6446000 ns,
x"01" after 6457000 ns,
x"93" after 6468000 ns,
x"F7" after 6479000 ns,
x"F7" after 6490000 ns,
x"0F" after 6501000 ns,
x"23" after 6512000 ns,
x"24" after 6523000 ns,
x"F4" after 6534000 ns,
x"FE" after 6545000 ns,
x"83" after 6556000 ns,
x"27" after 6567000 ns,
x"84" after 6578000 ns,
x"FE" after 6589000 ns,
x"63" after 6600000 ns,
x"88" after 6611000 ns,
x"07" after 6622000 ns,
x"00" after 6633000 ns,
x"83" after 6644000 ns,
x"27" after 6655000 ns,
x"04" after 6666000 ns,
x"FC" after 6677000 ns,
x"B3" after 6688000 ns,
x"07" after 6699000 ns,
x"F0" after 6710000 ns,
x"40" after 6721000 ns,
x"23" after 6732000 ns,
x"20" after 6743000 ns,
x"F4" after 6754000 ns,
x"FC" after 6765000 ns,
x"03" after 6776000 ns,
x"27" after 6787000 ns,
x"04" after 6798000 ns,
x"FC" after 6809000 ns,
x"93" after 6820000 ns,
x"07" after 6831000 ns,
x"A0" after 6842000 ns,
x"00" after 6853000 ns,
x"B3" after 6864000 ns,
x"67" after 6875000 ns,
x"F7" after 6886000 ns,
x"02" after 6897000 ns,
x"13" after 6908000 ns,
x"F7" after 6919000 ns,
x"F7" after 6930000 ns,
x"0F" after 6941000 ns,
x"83" after 6952000 ns,
x"27" after 6963000 ns,
x"44" after 6974000 ns,
x"FF" after 6985000 ns,
x"93" after 6996000 ns,
x"86" after 7007000 ns,
x"17" after 7018000 ns,
x"00" after 7029000 ns,
x"23" after 7040000 ns,
x"2A" after 7051000 ns,
x"D4" after 7062000 ns,
x"FE" after 7073000 ns,
x"13" after 7084000 ns,
x"07" after 7095000 ns,
x"07" after 7106000 ns,
x"03" after 7117000 ns,
x"13" after 7128000 ns,
x"77" after 7139000 ns,
x"F7" after 7150000 ns,
x"0F" after 7161000 ns,
x"93" after 7172000 ns,
x"87" after 7183000 ns,
x"87" after 7194000 ns,
x"FF" after 7205000 ns,
x"B3" after 7216000 ns,
x"87" after 7227000 ns,
x"87" after 7238000 ns,
x"00" after 7249000 ns,
x"23" after 7260000 ns,
x"88" after 7271000 ns,
x"E7" after 7282000 ns,
x"FC" after 7293000 ns,
x"03" after 7304000 ns,
x"27" after 7315000 ns,
x"04" after 7326000 ns,
x"FC" after 7337000 ns,
x"93" after 7348000 ns,
x"07" after 7359000 ns,
x"A0" after 7370000 ns,
x"00" after 7381000 ns,
x"B3" after 7392000 ns,
x"47" after 7403000 ns,
x"F7" after 7414000 ns,
x"02" after 7425000 ns,
x"23" after 7436000 ns,
x"20" after 7447000 ns,
x"F4" after 7458000 ns,
x"FC" after 7469000 ns,
x"83" after 7480000 ns,
x"27" after 7491000 ns,
x"04" after 7502000 ns,
x"FC" after 7513000 ns,
x"E3" after 7524000 ns,
x"9E" after 7535000 ns,
x"07" after 7546000 ns,
x"FA" after 7557000 ns,
x"83" after 7568000 ns,
x"27" after 7579000 ns,
x"84" after 7590000 ns,
x"FE" after 7601000 ns,
x"63" after 7612000 ns,
x"80" after 7623000 ns,
x"07" after 7634000 ns,
x"02" after 7645000 ns,
x"83" after 7656000 ns,
x"27" after 7667000 ns,
x"44" after 7678000 ns,
x"FF" after 7689000 ns,
x"13" after 7700000 ns,
x"87" after 7711000 ns,
x"17" after 7722000 ns,
x"00" after 7733000 ns,
x"23" after 7744000 ns,
x"2A" after 7755000 ns,
x"E4" after 7766000 ns,
x"FE" after 7777000 ns,
x"93" after 7788000 ns,
x"87" after 7799000 ns,
x"87" after 7810000 ns,
x"FF" after 7821000 ns,
x"B3" after 7832000 ns,
x"87" after 7843000 ns,
x"87" after 7854000 ns,
x"00" after 7865000 ns,
x"13" after 7876000 ns,
x"07" after 7887000 ns,
x"D0" after 7898000 ns,
x"02" after 7909000 ns,
x"23" after 7920000 ns,
x"88" after 7931000 ns,
x"E7" after 7942000 ns,
x"FC" after 7953000 ns,
x"83" after 7964000 ns,
x"27" after 7975000 ns,
x"44" after 7986000 ns,
x"FF" after 7997000 ns,
x"23" after 8008000 ns,
x"26" after 8019000 ns,
x"F4" after 8030000 ns,
x"FE" after 8041000 ns,
x"23" after 8052000 ns,
x"28" after 8063000 ns,
x"04" after 8074000 ns,
x"FE" after 8085000 ns,
x"6F" after 8096000 ns,
x"00" after 8107000 ns,
x"C0" after 8118000 ns,
x"03" after 8129000 ns,
x"83" after 8140000 ns,
x"27" after 8151000 ns,
x"C4" after 8162000 ns,
x"FE" after 8173000 ns,
x"13" after 8184000 ns,
x"87" after 8195000 ns,
x"F7" after 8206000 ns,
x"FF" after 8217000 ns,
x"83" after 8228000 ns,
x"27" after 8239000 ns,
x"04" after 8250000 ns,
x"FF" after 8261000 ns,
x"33" after 8272000 ns,
x"07" after 8283000 ns,
x"F7" after 8294000 ns,
x"40" after 8305000 ns,
x"83" after 8316000 ns,
x"27" after 8327000 ns,
x"04" after 8338000 ns,
x"FF" after 8349000 ns,
x"83" after 8360000 ns,
x"26" after 8371000 ns,
x"44" after 8382000 ns,
x"FC" after 8393000 ns,
x"B3" after 8404000 ns,
x"87" after 8415000 ns,
x"F6" after 8426000 ns,
x"00" after 8437000 ns,
x"13" after 8448000 ns,
x"07" after 8459000 ns,
x"87" after 8470000 ns,
x"FF" after 8481000 ns,
x"33" after 8492000 ns,
x"07" after 8503000 ns,
x"87" after 8514000 ns,
x"00" after 8525000 ns,
x"03" after 8536000 ns,
x"47" after 8547000 ns,
x"07" after 8558000 ns,
x"FD" after 8569000 ns,
x"23" after 8580000 ns,
x"80" after 8591000 ns,
x"E7" after 8602000 ns,
x"00" after 8613000 ns,
x"83" after 8624000 ns,
x"27" after 8635000 ns,
x"04" after 8646000 ns,
x"FF" after 8657000 ns,
x"93" after 8668000 ns,
x"87" after 8679000 ns,
x"17" after 8690000 ns,
x"00" after 8701000 ns,
x"23" after 8712000 ns,
x"28" after 8723000 ns,
x"F4" after 8734000 ns,
x"FE" after 8745000 ns,
x"03" after 8756000 ns,
x"27" after 8767000 ns,
x"04" after 8778000 ns,
x"FF" after 8789000 ns,
x"83" after 8800000 ns,
x"27" after 8811000 ns,
x"C4" after 8822000 ns,
x"FE" after 8833000 ns,
x"E3" after 8844000 ns,
x"40" after 8855000 ns,
x"F7" after 8866000 ns,
x"FC" after 8877000 ns,
x"83" after 8888000 ns,
x"27" after 8899000 ns,
x"C4" after 8910000 ns,
x"FE" after 8921000 ns,
x"03" after 8932000 ns,
x"27" after 8943000 ns,
x"44" after 8954000 ns,
x"FC" after 8965000 ns,
x"B3" after 8976000 ns,
x"07" after 8987000 ns,
x"F7" after 8998000 ns,
x"00" after 9009000 ns,
x"23" after 9020000 ns,
x"80" after 9031000 ns,
x"07" after 9042000 ns,
x"00" after 9053000 ns,
x"83" after 9064000 ns,
x"27" after 9075000 ns,
x"C4" after 9086000 ns,
x"FE" after 9097000 ns,
x"13" after 9108000 ns,
x"85" after 9119000 ns,
x"07" after 9130000 ns,
x"00" after 9141000 ns,
x"03" after 9152000 ns,
x"24" after 9163000 ns,
x"C1" after 9174000 ns,
x"03" after 9185000 ns,
x"13" after 9196000 ns,
x"01" after 9207000 ns,
x"01" after 9218000 ns,
x"04" after 9229000 ns,
x"67" after 9240000 ns,
x"80" after 9251000 ns,
x"00" after 9262000 ns,
x"00" after 9273000 ns,
x"13" after 9284000 ns,
x"01" after 9295000 ns,
x"01" after 9306000 ns,
x"FB" after 9317000 ns,
x"23" after 9328000 ns,
x"2A" after 9339000 ns,
x"11" after 9350000 ns,
x"02" after 9361000 ns,
x"23" after 9372000 ns,
x"28" after 9383000 ns,
x"81" after 9394000 ns,
x"02" after 9405000 ns,
x"13" after 9416000 ns,
x"04" after 9427000 ns,
x"81" after 9438000 ns,
x"03" after 9449000 ns,
x"23" after 9460000 ns,
x"2A" after 9471000 ns,
x"A4" after 9482000 ns,
x"FC" after 9493000 ns,
x"23" after 9504000 ns,
x"28" after 9515000 ns,
x"B4" after 9526000 ns,
x"FC" after 9537000 ns,
x"23" after 9548000 ns,
x"20" after 9559000 ns,
x"C4" after 9570000 ns,
x"00" after 9581000 ns,
x"23" after 9592000 ns,
x"22" after 9603000 ns,
x"D4" after 9614000 ns,
x"00" after 9625000 ns,
x"23" after 9636000 ns,
x"24" after 9647000 ns,
x"E4" after 9658000 ns,
x"00" after 9669000 ns,
x"23" after 9680000 ns,
x"26" after 9691000 ns,
x"F4" after 9702000 ns,
x"00" after 9713000 ns,
x"23" after 9724000 ns,
x"28" after 9735000 ns,
x"04" after 9746000 ns,
x"01" after 9757000 ns,
x"23" after 9768000 ns,
x"2A" after 9779000 ns,
x"14" after 9790000 ns,
x"01" after 9801000 ns,
x"93" after 9812000 ns,
x"07" after 9823000 ns,
x"84" after 9834000 ns,
x"01" after 9845000 ns,
x"23" after 9856000 ns,
x"26" after 9867000 ns,
x"F4" after 9878000 ns,
x"FC" after 9889000 ns,
x"83" after 9900000 ns,
x"27" after 9911000 ns,
x"C4" after 9922000 ns,
x"FC" after 9933000 ns,
x"93" after 9944000 ns,
x"87" after 9955000 ns,
x"87" after 9966000 ns,
x"FE" after 9977000 ns,
x"23" after 9988000 ns,
x"2E" after 9999000 ns,
x"F4" after 10010000 ns,
x"FC" after 10021000 ns,
x"83" after 10032000 ns,
x"27" after 10043000 ns,
x"04" after 10054000 ns,
x"FD" after 10065000 ns,
x"23" after 10076000 ns,
x"2A" after 10087000 ns,
x"F4" after 10098000 ns,
x"FE" after 10109000 ns,
x"83" after 10120000 ns,
x"27" after 10131000 ns,
x"44" after 10142000 ns,
x"FD" after 10153000 ns,
x"23" after 10164000 ns,
x"28" after 10175000 ns,
x"F4" after 10186000 ns,
x"FE" after 10197000 ns,
x"6F" after 10208000 ns,
x"00" after 10219000 ns,
x"00" after 10230000 ns,
x"21" after 10241000 ns,
x"83" after 10252000 ns,
x"27" after 10263000 ns,
x"44" after 10274000 ns,
x"FF" after 10285000 ns,
x"03" after 10296000 ns,
x"C7" after 10307000 ns,
x"07" after 10318000 ns,
x"00" after 10329000 ns,
x"93" after 10340000 ns,
x"07" after 10351000 ns,
x"50" after 10362000 ns,
x"02" after 10373000 ns,
x"63" after 10384000 ns,
x"1E" after 10395000 ns,
x"F7" after 10406000 ns,
x"1C" after 10417000 ns,
x"83" after 10428000 ns,
x"27" after 10439000 ns,
x"44" after 10450000 ns,
x"FF" after 10461000 ns,
x"93" after 10472000 ns,
x"87" after 10483000 ns,
x"17" after 10494000 ns,
x"00" after 10505000 ns,
x"23" after 10516000 ns,
x"2A" after 10527000 ns,
x"F4" after 10538000 ns,
x"FE" after 10549000 ns,
x"83" after 10560000 ns,
x"27" after 10571000 ns,
x"44" after 10582000 ns,
x"FF" after 10593000 ns,
x"83" after 10604000 ns,
x"C7" after 10615000 ns,
x"07" after 10626000 ns,
x"00" after 10637000 ns,
x"13" after 10648000 ns,
x"07" after 10659000 ns,
x"30" after 10670000 ns,
x"07" after 10681000 ns,
x"63" after 10692000 ns,
x"8C" after 10703000 ns,
x"E7" after 10714000 ns,
x"06" after 10725000 ns,
x"13" after 10736000 ns,
x"07" after 10747000 ns,
x"30" after 10758000 ns,
x"07" after 10769000 ns,
x"63" after 10780000 ns,
x"44" after 10791000 ns,
x"F7" after 10802000 ns,
x"18" after 10813000 ns,
x"13" after 10824000 ns,
x"07" after 10835000 ns,
x"40" after 10846000 ns,
x"06" after 10857000 ns,
x"63" after 10868000 ns,
x"88" after 10879000 ns,
x"E7" after 10890000 ns,
x"02" after 10901000 ns,
x"13" after 10912000 ns,
x"07" after 10923000 ns,
x"40" after 10934000 ns,
x"06" after 10945000 ns,
x"63" after 10956000 ns,
x"4C" after 10967000 ns,
x"F7" after 10978000 ns,
x"16" after 10989000 ns,
x"13" after 11000000 ns,
x"07" after 11011000 ns,
x"30" after 11022000 ns,
x"06" after 11033000 ns,
x"63" after 11044000 ns,
x"88" after 11055000 ns,
x"E7" after 11066000 ns,
x"08" after 11077000 ns,
x"13" after 11088000 ns,
x"07" after 11099000 ns,
x"30" after 11110000 ns,
x"06" after 11121000 ns,
x"63" after 11132000 ns,
x"44" after 11143000 ns,
x"F7" after 11154000 ns,
x"16" after 11165000 ns,
x"13" after 11176000 ns,
x"07" after 11187000 ns,
x"50" after 11198000 ns,
x"02" after 11209000 ns,
x"63" after 11220000 ns,
x"86" after 11231000 ns,
x"E7" after 11242000 ns,
x"0A" after 11253000 ns,
x"13" after 11264000 ns,
x"07" after 11275000 ns,
x"00" after 11286000 ns,
x"03" after 11297000 ns,
x"63" after 11308000 ns,
x"8E" after 11319000 ns,
x"E7" after 11330000 ns,
x"0A" after 11341000 ns,
x"6F" after 11352000 ns,
x"00" after 11363000 ns,
x"40" after 11374000 ns,
x"15" after 11385000 ns,
x"83" after 11396000 ns,
x"27" after 11407000 ns,
x"C4" after 11418000 ns,
x"FD" after 11429000 ns,
x"13" after 11440000 ns,
x"87" after 11451000 ns,
x"47" after 11462000 ns,
x"00" after 11473000 ns,
x"23" after 11484000 ns,
x"2E" after 11495000 ns,
x"E4" after 11506000 ns,
x"FC" after 11517000 ns,
x"83" after 11528000 ns,
x"A7" after 11539000 ns,
x"07" after 11550000 ns,
x"00" after 11561000 ns,
x"23" after 11572000 ns,
x"24" after 11583000 ns,
x"F4" after 11594000 ns,
x"FE" after 11605000 ns,
x"83" after 11616000 ns,
x"25" after 11627000 ns,
x"84" after 11638000 ns,
x"FE" after 11649000 ns,
x"03" after 11660000 ns,
x"25" after 11671000 ns,
x"04" after 11682000 ns,
x"FF" after 11693000 ns,
x"EF" after 11704000 ns,
x"F0" after 11715000 ns,
x"1F" after 11726000 ns,
x"E0" after 11737000 ns,
x"93" after 11748000 ns,
x"07" after 11759000 ns,
x"05" after 11770000 ns,
x"00" after 11781000 ns,
x"13" after 11792000 ns,
x"87" after 11803000 ns,
x"07" after 11814000 ns,
x"00" after 11825000 ns,
x"83" after 11836000 ns,
x"27" after 11847000 ns,
x"04" after 11858000 ns,
x"FF" after 11869000 ns,
x"B3" after 11880000 ns,
x"87" after 11891000 ns,
x"E7" after 11902000 ns,
x"00" after 11913000 ns,
x"23" after 11924000 ns,
x"28" after 11935000 ns,
x"F4" after 11946000 ns,
x"FE" after 11957000 ns,
x"6F" after 11968000 ns,
x"00" after 11979000 ns,
x"40" after 11990000 ns,
x"16" after 12001000 ns,
x"83" after 12012000 ns,
x"27" after 12023000 ns,
x"C4" after 12034000 ns,
x"FD" after 12045000 ns,
x"13" after 12056000 ns,
x"87" after 12067000 ns,
x"47" after 12078000 ns,
x"00" after 12089000 ns,
x"23" after 12100000 ns,
x"2E" after 12111000 ns,
x"E4" after 12122000 ns,
x"FC" after 12133000 ns,
x"83" after 12144000 ns,
x"A7" after 12155000 ns,
x"07" after 12166000 ns,
x"00" after 12177000 ns,
x"23" after 12188000 ns,
x"26" after 12199000 ns,
x"F4" after 12210000 ns,
x"FE" after 12221000 ns,
x"83" after 12232000 ns,
x"25" after 12243000 ns,
x"C4" after 12254000 ns,
x"FE" after 12265000 ns,
x"03" after 12276000 ns,
x"25" after 12287000 ns,
x"04" after 12298000 ns,
x"FF" after 12309000 ns,
x"EF" after 12320000 ns,
x"F0" after 12331000 ns,
x"5F" after 12342000 ns,
x"CB" after 12353000 ns,
x"93" after 12364000 ns,
x"07" after 12375000 ns,
x"05" after 12386000 ns,
x"00" after 12397000 ns,
x"13" after 12408000 ns,
x"87" after 12419000 ns,
x"07" after 12430000 ns,
x"00" after 12441000 ns,
x"83" after 12452000 ns,
x"27" after 12463000 ns,
x"04" after 12474000 ns,
x"FF" after 12485000 ns,
x"B3" after 12496000 ns,
x"87" after 12507000 ns,
x"E7" after 12518000 ns,
x"00" after 12529000 ns,
x"23" after 12540000 ns,
x"28" after 12551000 ns,
x"F4" after 12562000 ns,
x"FE" after 12573000 ns,
x"6F" after 12584000 ns,
x"00" after 12595000 ns,
x"C0" after 12606000 ns,
x"12" after 12617000 ns,
x"83" after 12628000 ns,
x"27" after 12639000 ns,
x"C4" after 12650000 ns,
x"FD" after 12661000 ns,
x"13" after 12672000 ns,
x"87" after 12683000 ns,
x"47" after 12694000 ns,
x"00" after 12705000 ns,
x"23" after 12716000 ns,
x"2E" after 12727000 ns,
x"E4" after 12738000 ns,
x"FC" after 12749000 ns,
x"83" after 12760000 ns,
x"A7" after 12771000 ns,
x"07" after 12782000 ns,
x"00" after 12793000 ns,
x"A3" after 12804000 ns,
x"03" after 12815000 ns,
x"F4" after 12826000 ns,
x"FE" after 12837000 ns,
x"83" after 12848000 ns,
x"27" after 12859000 ns,
x"04" after 12870000 ns,
x"FF" after 12881000 ns,
x"13" after 12892000 ns,
x"87" after 12903000 ns,
x"17" after 12914000 ns,
x"00" after 12925000 ns,
x"23" after 12936000 ns,
x"28" after 12947000 ns,
x"E4" after 12958000 ns,
x"FE" after 12969000 ns,
x"03" after 12980000 ns,
x"47" after 12991000 ns,
x"74" after 13002000 ns,
x"FE" after 13013000 ns,
x"23" after 13024000 ns,
x"80" after 13035000 ns,
x"E7" after 13046000 ns,
x"00" after 13057000 ns,
x"6F" after 13068000 ns,
x"00" after 13079000 ns,
x"00" after 13090000 ns,
x"10" after 13101000 ns,
x"83" after 13112000 ns,
x"27" after 13123000 ns,
x"04" after 13134000 ns,
x"FF" after 13145000 ns,
x"13" after 13156000 ns,
x"87" after 13167000 ns,
x"17" after 13178000 ns,
x"00" after 13189000 ns,
x"23" after 13200000 ns,
x"28" after 13211000 ns,
x"E4" after 13222000 ns,
x"FE" after 13233000 ns,
x"13" after 13244000 ns,
x"07" after 13255000 ns,
x"50" after 13266000 ns,
x"02" after 13277000 ns,
x"23" after 13288000 ns,
x"80" after 13299000 ns,
x"E7" after 13310000 ns,
x"00" after 13321000 ns,
x"6F" after 13332000 ns,
x"00" after 13343000 ns,
x"80" after 13354000 ns,
x"0E" after 13365000 ns,
x"83" after 13376000 ns,
x"27" after 13387000 ns,
x"44" after 13398000 ns,
x"FF" after 13409000 ns,
x"93" after 13420000 ns,
x"87" after 13431000 ns,
x"17" after 13442000 ns,
x"00" after 13453000 ns,
x"03" after 13464000 ns,
x"C7" after 13475000 ns,
x"07" after 13486000 ns,
x"00" after 13497000 ns,
x"93" after 13508000 ns,
x"07" after 13519000 ns,
x"20" after 13530000 ns,
x"03" after 13541000 ns,
x"63" after 13552000 ns,
x"10" after 13563000 ns,
x"F7" after 13574000 ns,
x"06" after 13585000 ns,
x"83" after 13596000 ns,
x"27" after 13607000 ns,
x"44" after 13618000 ns,
x"FF" after 13629000 ns,
x"93" after 13640000 ns,
x"87" after 13651000 ns,
x"27" after 13662000 ns,
x"00" after 13673000 ns,
x"03" after 13684000 ns,
x"C7" after 13695000 ns,
x"07" after 13706000 ns,
x"00" after 13717000 ns,
x"93" after 13728000 ns,
x"07" after 13739000 ns,
x"80" after 13750000 ns,
x"05" after 13761000 ns,
x"63" after 13772000 ns,
x"16" after 13783000 ns,
x"F7" after 13794000 ns,
x"04" after 13805000 ns,
x"83" after 13816000 ns,
x"27" after 13827000 ns,
x"44" after 13838000 ns,
x"FF" after 13849000 ns,
x"93" after 13860000 ns,
x"87" after 13871000 ns,
x"27" after 13882000 ns,
x"00" after 13893000 ns,
x"23" after 13904000 ns,
x"2A" after 13915000 ns,
x"F4" after 13926000 ns,
x"FE" after 13937000 ns,
x"83" after 13948000 ns,
x"27" after 13959000 ns,
x"C4" after 13970000 ns,
x"FD" after 13981000 ns,
x"13" after 13992000 ns,
x"87" after 14003000 ns,
x"47" after 14014000 ns,
x"00" after 14025000 ns,
x"23" after 14036000 ns,
x"2E" after 14047000 ns,
x"E4" after 14058000 ns,
x"FC" after 14069000 ns,
x"83" after 14080000 ns,
x"A7" after 14091000 ns,
x"07" after 14102000 ns,
x"00" after 14113000 ns,
x"23" after 14124000 ns,
x"20" after 14135000 ns,
x"F4" after 14146000 ns,
x"FE" after 14157000 ns,
x"83" after 14168000 ns,
x"25" after 14179000 ns,
x"04" after 14190000 ns,
x"FE" after 14201000 ns,
x"03" after 14212000 ns,
x"25" after 14223000 ns,
x"04" after 14234000 ns,
x"FF" after 14245000 ns,
x"EF" after 14256000 ns,
x"F0" after 14267000 ns,
x"5F" after 14278000 ns,
x"C7" after 14289000 ns,
x"93" after 14300000 ns,
x"07" after 14311000 ns,
x"05" after 14322000 ns,
x"00" after 14333000 ns,
x"13" after 14344000 ns,
x"87" after 14355000 ns,
x"07" after 14366000 ns,
x"00" after 14377000 ns,
x"83" after 14388000 ns,
x"27" after 14399000 ns,
x"04" after 14410000 ns,
x"FF" after 14421000 ns,
x"B3" after 14432000 ns,
x"87" after 14443000 ns,
x"E7" after 14454000 ns,
x"00" after 14465000 ns,
x"23" after 14476000 ns,
x"28" after 14487000 ns,
x"F4" after 14498000 ns,
x"FE" after 14509000 ns,
x"13" after 14520000 ns,
x"00" after 14531000 ns,
x"00" after 14542000 ns,
x"00" after 14553000 ns,
x"6F" after 14564000 ns,
x"00" after 14575000 ns,
x"80" after 14586000 ns,
x"07" after 14597000 ns,
x"83" after 14608000 ns,
x"27" after 14619000 ns,
x"04" after 14630000 ns,
x"FF" after 14641000 ns,
x"13" after 14652000 ns,
x"87" after 14663000 ns,
x"17" after 14674000 ns,
x"00" after 14685000 ns,
x"23" after 14696000 ns,
x"28" after 14707000 ns,
x"E4" after 14718000 ns,
x"FE" after 14729000 ns,
x"13" after 14740000 ns,
x"07" after 14751000 ns,
x"50" after 14762000 ns,
x"02" after 14773000 ns,
x"23" after 14784000 ns,
x"80" after 14795000 ns,
x"E7" after 14806000 ns,
x"00" after 14817000 ns,
x"83" after 14828000 ns,
x"27" after 14839000 ns,
x"04" after 14850000 ns,
x"FF" after 14861000 ns,
x"13" after 14872000 ns,
x"87" after 14883000 ns,
x"17" after 14894000 ns,
x"00" after 14905000 ns,
x"23" after 14916000 ns,
x"28" after 14927000 ns,
x"E4" after 14938000 ns,
x"FE" after 14949000 ns,
x"13" after 14960000 ns,
x"07" after 14971000 ns,
x"00" after 14982000 ns,
x"03" after 14993000 ns,
x"23" after 15004000 ns,
x"80" after 15015000 ns,
x"E7" after 15026000 ns,
x"00" after 15037000 ns,
x"6F" after 15048000 ns,
x"00" after 15059000 ns,
x"C0" after 15070000 ns,
x"04" after 15081000 ns,
x"83" after 15092000 ns,
x"27" after 15103000 ns,
x"04" after 15114000 ns,
x"FF" after 15125000 ns,
x"13" after 15136000 ns,
x"87" after 15147000 ns,
x"17" after 15158000 ns,
x"00" after 15169000 ns,
x"23" after 15180000 ns,
x"28" after 15191000 ns,
x"E4" after 15202000 ns,
x"FE" after 15213000 ns,
x"13" after 15224000 ns,
x"07" after 15235000 ns,
x"50" after 15246000 ns,
x"02" after 15257000 ns,
x"23" after 15268000 ns,
x"80" after 15279000 ns,
x"E7" after 15290000 ns,
x"00" after 15301000 ns,
x"83" after 15312000 ns,
x"27" after 15323000 ns,
x"04" after 15334000 ns,
x"FF" after 15345000 ns,
x"13" after 15356000 ns,
x"87" after 15367000 ns,
x"17" after 15378000 ns,
x"00" after 15389000 ns,
x"23" after 15400000 ns,
x"28" after 15411000 ns,
x"E4" after 15422000 ns,
x"FE" after 15433000 ns,
x"03" after 15444000 ns,
x"27" after 15455000 ns,
x"44" after 15466000 ns,
x"FF" after 15477000 ns,
x"03" after 15488000 ns,
x"47" after 15499000 ns,
x"07" after 15510000 ns,
x"00" after 15521000 ns,
x"23" after 15532000 ns,
x"80" after 15543000 ns,
x"E7" after 15554000 ns,
x"00" after 15565000 ns,
x"6F" after 15576000 ns,
x"00" after 15587000 ns,
x"C0" after 15598000 ns,
x"01" after 15609000 ns,
x"83" after 15620000 ns,
x"27" after 15631000 ns,
x"04" after 15642000 ns,
x"FF" after 15653000 ns,
x"13" after 15664000 ns,
x"87" after 15675000 ns,
x"17" after 15686000 ns,
x"00" after 15697000 ns,
x"23" after 15708000 ns,
x"28" after 15719000 ns,
x"E4" after 15730000 ns,
x"FE" after 15741000 ns,
x"03" after 15752000 ns,
x"27" after 15763000 ns,
x"44" after 15774000 ns,
x"FF" after 15785000 ns,
x"03" after 15796000 ns,
x"47" after 15807000 ns,
x"07" after 15818000 ns,
x"00" after 15829000 ns,
x"23" after 15840000 ns,
x"80" after 15851000 ns,
x"E7" after 15862000 ns,
x"00" after 15873000 ns,
x"83" after 15884000 ns,
x"27" after 15895000 ns,
x"44" after 15906000 ns,
x"FF" after 15917000 ns,
x"93" after 15928000 ns,
x"87" after 15939000 ns,
x"17" after 15950000 ns,
x"00" after 15961000 ns,
x"23" after 15972000 ns,
x"2A" after 15983000 ns,
x"F4" after 15994000 ns,
x"FE" after 16005000 ns,
x"83" after 16016000 ns,
x"27" after 16027000 ns,
x"44" after 16038000 ns,
x"FF" after 16049000 ns,
x"83" after 16060000 ns,
x"C7" after 16071000 ns,
x"07" after 16082000 ns,
x"00" after 16093000 ns,
x"E3" after 16104000 ns,
x"96" after 16115000 ns,
x"07" after 16126000 ns,
x"DE" after 16137000 ns,
x"83" after 16148000 ns,
x"27" after 16159000 ns,
x"04" after 16170000 ns,
x"FF" after 16181000 ns,
x"23" after 16192000 ns,
x"80" after 16203000 ns,
x"07" after 16214000 ns,
x"00" after 16225000 ns,
x"13" after 16236000 ns,
x"00" after 16247000 ns,
x"00" after 16258000 ns,
x"00" after 16269000 ns,
x"83" after 16280000 ns,
x"20" after 16291000 ns,
x"41" after 16302000 ns,
x"03" after 16313000 ns,
x"03" after 16324000 ns,
x"24" after 16335000 ns,
x"01" after 16346000 ns,
x"03" after 16357000 ns,
x"13" after 16368000 ns,
x"01" after 16379000 ns,
x"01" after 16390000 ns,
x"05" after 16401000 ns,
x"67" after 16412000 ns,
x"80" after 16423000 ns,
x"00" after 16434000 ns,
x"00" after 16445000 ns,
x"13" after 16456000 ns,
x"01" after 16467000 ns,
x"01" after 16478000 ns,
x"FF" after 16489000 ns,
x"23" after 16500000 ns,
x"26" after 16511000 ns,
x"81" after 16522000 ns,
x"00" after 16533000 ns,
x"13" after 16544000 ns,
x"04" after 16555000 ns,
x"01" after 16566000 ns,
x"01" after 16577000 ns,
x"23" after 16588000 ns,
x"2A" after 16599000 ns,
x"A4" after 16610000 ns,
x"FE" after 16621000 ns,
x"6F" after 16632000 ns,
x"00" after 16643000 ns,
x"00" after 16654000 ns,
x"01" after 16665000 ns,
x"83" after 16676000 ns,
x"27" after 16687000 ns,
x"44" after 16698000 ns,
x"FF" after 16709000 ns,
x"93" after 16720000 ns,
x"87" after 16731000 ns,
x"F7" after 16742000 ns,
x"FF" after 16753000 ns,
x"23" after 16764000 ns,
x"2A" after 16775000 ns,
x"F4" after 16786000 ns,
x"FE" after 16797000 ns,
x"83" after 16808000 ns,
x"27" after 16819000 ns,
x"44" after 16830000 ns,
x"FF" after 16841000 ns,
x"E3" after 16852000 ns,
x"48" after 16863000 ns,
x"F0" after 16874000 ns,
x"FE" after 16885000 ns,
x"13" after 16896000 ns,
x"00" after 16907000 ns,
x"00" after 16918000 ns,
x"00" after 16929000 ns,
x"13" after 16940000 ns,
x"00" after 16951000 ns,
x"00" after 16962000 ns,
x"00" after 16973000 ns,
x"03" after 16984000 ns,
x"24" after 16995000 ns,
x"C1" after 17006000 ns,
x"00" after 17017000 ns,
x"13" after 17028000 ns,
x"01" after 17039000 ns,
x"01" after 17050000 ns,
x"01" after 17061000 ns,
x"67" after 17072000 ns,
x"80" after 17083000 ns,
x"00" after 17094000 ns,
x"00" after 17105000 ns,
x"13" after 17116000 ns,
x"01" after 17127000 ns,
x"01" after 17138000 ns,
x"FF" after 17149000 ns,
x"23" after 17160000 ns,
x"26" after 17171000 ns,
x"11" after 17182000 ns,
x"00" after 17193000 ns,
x"23" after 17204000 ns,
x"24" after 17215000 ns,
x"81" after 17226000 ns,
x"00" after 17237000 ns,
x"13" after 17248000 ns,
x"04" after 17259000 ns,
x"01" after 17270000 ns,
x"01" after 17281000 ns,
x"B7" after 17292000 ns,
x"17" after 17303000 ns,
x"00" after 17314000 ns,
x"00" after 17325000 ns,
x"93" after 17336000 ns,
x"87" after 17347000 ns,
x"07" after 17358000 ns,
x"80" after 17369000 ns,
x"83" after 17380000 ns,
x"A7" after 17391000 ns,
x"07" after 17402000 ns,
x"00" after 17413000 ns,
x"37" after 17424000 ns,
x"17" after 17435000 ns,
x"00" after 17446000 ns,
x"00" after 17457000 ns,
x"13" after 17468000 ns,
x"07" after 17479000 ns,
x"07" after 17490000 ns,
x"81" after 17501000 ns,
x"93" after 17512000 ns,
x"97" after 17523000 ns,
x"27" after 17534000 ns,
x"00" after 17545000 ns,
x"B3" after 17556000 ns,
x"07" after 17567000 ns,
x"F7" after 17578000 ns,
x"00" after 17589000 ns,
x"83" after 17600000 ns,
x"A7" after 17611000 ns,
x"07" after 17622000 ns,
x"00" after 17633000 ns,
x"23" after 17644000 ns,
x"2A" after 17655000 ns,
x"F4" after 17666000 ns,
x"FE" after 17677000 ns,
x"83" after 17688000 ns,
x"27" after 17699000 ns,
x"44" after 17710000 ns,
x"FF" after 17721000 ns,
x"93" after 17732000 ns,
x"E7" after 17743000 ns,
x"77" after 17754000 ns,
x"00" after 17765000 ns,
x"23" after 17776000 ns,
x"2A" after 17787000 ns,
x"F4" after 17798000 ns,
x"FE" after 17809000 ns,
x"03" after 17820000 ns,
x"25" after 17831000 ns,
x"44" after 17842000 ns,
x"FF" after 17853000 ns,
x"EF" after 17864000 ns,
x"F0" after 17875000 ns,
x"1F" after 17886000 ns,
x"A3" after 17897000 ns,
x"B7" after 17908000 ns,
x"67" after 17919000 ns,
x"00" after 17930000 ns,
x"00" after 17941000 ns,
x"13" after 17952000 ns,
x"85" after 17963000 ns,
x"87" after 17974000 ns,
x"1A" after 17985000 ns,
x"EF" after 17996000 ns,
x"F0" after 18007000 ns,
x"5F" after 18018000 ns,
x"F7" after 18029000 ns,
x"B7" after 18040000 ns,
x"17" after 18051000 ns,
x"00" after 18062000 ns,
x"00" after 18073000 ns,
x"93" after 18084000 ns,
x"87" after 18095000 ns,
x"07" after 18106000 ns,
x"80" after 18117000 ns,
x"83" after 18128000 ns,
x"A7" after 18139000 ns,
x"47" after 18150000 ns,
x"00" after 18161000 ns,
x"37" after 18172000 ns,
x"17" after 18183000 ns,
x"00" after 18194000 ns,
x"00" after 18205000 ns,
x"13" after 18216000 ns,
x"07" after 18227000 ns,
x"07" after 18238000 ns,
x"81" after 18249000 ns,
x"93" after 18260000 ns,
x"97" after 18271000 ns,
x"27" after 18282000 ns,
x"00" after 18293000 ns,
x"B3" after 18304000 ns,
x"07" after 18315000 ns,
x"F7" after 18326000 ns,
x"00" after 18337000 ns,
x"83" after 18348000 ns,
x"A7" after 18359000 ns,
x"07" after 18370000 ns,
x"00" after 18381000 ns,
x"23" after 18392000 ns,
x"2A" after 18403000 ns,
x"F4" after 18414000 ns,
x"FE" after 18425000 ns,
x"83" after 18436000 ns,
x"27" after 18447000 ns,
x"44" after 18458000 ns,
x"FF" after 18469000 ns,
x"93" after 18480000 ns,
x"E7" after 18491000 ns,
x"B7" after 18502000 ns,
x"00" after 18513000 ns,
x"23" after 18524000 ns,
x"2A" after 18535000 ns,
x"F4" after 18546000 ns,
x"FE" after 18557000 ns,
x"03" after 18568000 ns,
x"25" after 18579000 ns,
x"44" after 18590000 ns,
x"FF" after 18601000 ns,
x"EF" after 18612000 ns,
x"F0" after 18623000 ns,
x"DF" after 18634000 ns,
x"9E" after 18645000 ns,
x"B7" after 18656000 ns,
x"67" after 18667000 ns,
x"00" after 18678000 ns,
x"00" after 18689000 ns,
x"13" after 18700000 ns,
x"85" after 18711000 ns,
x"87" after 18722000 ns,
x"1A" after 18733000 ns,
x"EF" after 18744000 ns,
x"F0" after 18755000 ns,
x"1F" after 18766000 ns,
x"F3" after 18777000 ns,
x"B7" after 18788000 ns,
x"17" after 18799000 ns,
x"00" after 18810000 ns,
x"00" after 18821000 ns,
x"93" after 18832000 ns,
x"87" after 18843000 ns,
x"07" after 18854000 ns,
x"80" after 18865000 ns,
x"83" after 18876000 ns,
x"A7" after 18887000 ns,
x"87" after 18898000 ns,
x"00" after 18909000 ns,
x"37" after 18920000 ns,
x"17" after 18931000 ns,
x"00" after 18942000 ns,
x"00" after 18953000 ns,
x"13" after 18964000 ns,
x"07" after 18975000 ns,
x"07" after 18986000 ns,
x"81" after 18997000 ns,
x"93" after 19008000 ns,
x"97" after 19019000 ns,
x"27" after 19030000 ns,
x"00" after 19041000 ns,
x"B3" after 19052000 ns,
x"07" after 19063000 ns,
x"F7" after 19074000 ns,
x"00" after 19085000 ns,
x"83" after 19096000 ns,
x"A7" after 19107000 ns,
x"07" after 19118000 ns,
x"00" after 19129000 ns,
x"23" after 19140000 ns,
x"2A" after 19151000 ns,
x"F4" after 19162000 ns,
x"FE" after 19173000 ns,
x"83" after 19184000 ns,
x"27" after 19195000 ns,
x"44" after 19206000 ns,
x"FF" after 19217000 ns,
x"93" after 19228000 ns,
x"E7" after 19239000 ns,
x"D7" after 19250000 ns,
x"00" after 19261000 ns,
x"23" after 19272000 ns,
x"2A" after 19283000 ns,
x"F4" after 19294000 ns,
x"FE" after 19305000 ns,
x"03" after 19316000 ns,
x"25" after 19327000 ns,
x"44" after 19338000 ns,
x"FF" after 19349000 ns,
x"EF" after 19360000 ns,
x"F0" after 19371000 ns,
x"9F" after 19382000 ns,
x"9A" after 19393000 ns,
x"B7" after 19404000 ns,
x"67" after 19415000 ns,
x"00" after 19426000 ns,
x"00" after 19437000 ns,
x"13" after 19448000 ns,
x"85" after 19459000 ns,
x"87" after 19470000 ns,
x"1A" after 19481000 ns,
x"EF" after 19492000 ns,
x"F0" after 19503000 ns,
x"DF" after 19514000 ns,
x"EE" after 19525000 ns,
x"B7" after 19536000 ns,
x"17" after 19547000 ns,
x"00" after 19558000 ns,
x"00" after 19569000 ns,
x"93" after 19580000 ns,
x"87" after 19591000 ns,
x"07" after 19602000 ns,
x"80" after 19613000 ns,
x"83" after 19624000 ns,
x"A7" after 19635000 ns,
x"C7" after 19646000 ns,
x"00" after 19657000 ns,
x"37" after 19668000 ns,
x"17" after 19679000 ns,
x"00" after 19690000 ns,
x"00" after 19701000 ns,
x"13" after 19712000 ns,
x"07" after 19723000 ns,
x"07" after 19734000 ns,
x"81" after 19745000 ns,
x"93" after 19756000 ns,
x"97" after 19767000 ns,
x"27" after 19778000 ns,
x"00" after 19789000 ns,
x"B3" after 19800000 ns,
x"07" after 19811000 ns,
x"F7" after 19822000 ns,
x"00" after 19833000 ns,
x"83" after 19844000 ns,
x"A7" after 19855000 ns,
x"07" after 19866000 ns,
x"00" after 19877000 ns,
x"23" after 19888000 ns,
x"2A" after 19899000 ns,
x"F4" after 19910000 ns,
x"FE" after 19921000 ns,
x"83" after 19932000 ns,
x"27" after 19943000 ns,
x"44" after 19954000 ns,
x"FF" after 19965000 ns,
x"93" after 19976000 ns,
x"E7" after 19987000 ns,
x"E7" after 19998000 ns,
x"00" after 20009000 ns,
x"23" after 20020000 ns,
x"2A" after 20031000 ns,
x"F4" after 20042000 ns,
x"FE" after 20053000 ns,
x"03" after 20064000 ns,
x"25" after 20075000 ns,
x"44" after 20086000 ns,
x"FF" after 20097000 ns,
x"EF" after 20108000 ns,
x"F0" after 20119000 ns,
x"5F" after 20130000 ns,
x"96" after 20141000 ns,
x"13" after 20152000 ns,
x"00" after 20163000 ns,
x"00" after 20174000 ns,
x"00" after 20185000 ns,
x"83" after 20196000 ns,
x"20" after 20207000 ns,
x"C1" after 20218000 ns,
x"00" after 20229000 ns,
x"03" after 20240000 ns,
x"24" after 20251000 ns,
x"81" after 20262000 ns,
x"00" after 20273000 ns,
x"13" after 20284000 ns,
x"01" after 20295000 ns,
x"01" after 20306000 ns,
x"01" after 20317000 ns,
x"67" after 20328000 ns,
x"80" after 20339000 ns,
x"00" after 20350000 ns,
x"00" after 20361000 ns,
x"13" after 20372000 ns,
x"01" after 20383000 ns,
x"01" after 20394000 ns,
x"FF" after 20405000 ns,
x"23" after 20416000 ns,
x"26" after 20427000 ns,
x"81" after 20438000 ns,
x"00" after 20449000 ns,
x"13" after 20460000 ns,
x"04" after 20471000 ns,
x"01" after 20482000 ns,
x"01" after 20493000 ns,
x"23" after 20504000 ns,
x"2A" after 20515000 ns,
x"04" after 20526000 ns,
x"FE" after 20537000 ns,
x"6F" after 20548000 ns,
x"00" after 20559000 ns,
x"00" after 20570000 ns,
x"01" after 20581000 ns,
x"83" after 20592000 ns,
x"27" after 20603000 ns,
x"44" after 20614000 ns,
x"FF" after 20625000 ns,
x"93" after 20636000 ns,
x"87" after 20647000 ns,
x"17" after 20658000 ns,
x"00" after 20669000 ns,
x"23" after 20680000 ns,
x"2A" after 20691000 ns,
x"F4" after 20702000 ns,
x"FE" after 20713000 ns,
x"03" after 20724000 ns,
x"27" after 20735000 ns,
x"44" after 20746000 ns,
x"FF" after 20757000 ns,
x"B7" after 20768000 ns,
x"C7" after 20779000 ns,
x"0D" after 20790000 ns,
x"00" after 20801000 ns,
x"93" after 20812000 ns,
x"87" after 20823000 ns,
x"F7" after 20834000 ns,
x"B9" after 20845000 ns,
x"E3" after 20856000 ns,
x"D4" after 20867000 ns,
x"E7" after 20878000 ns,
x"FE" after 20889000 ns,
x"B7" after 20900000 ns,
x"17" after 20911000 ns,
x"00" after 20922000 ns,
x"00" after 20933000 ns,
x"83" after 20944000 ns,
x"A7" after 20955000 ns,
x"47" after 20966000 ns,
x"85" after 20977000 ns,
x"13" after 20988000 ns,
x"87" after 20999000 ns,
x"F7" after 21010000 ns,
x"FF" after 21021000 ns,
x"B7" after 21032000 ns,
x"17" after 21043000 ns,
x"00" after 21054000 ns,
x"00" after 21065000 ns,
x"23" after 21076000 ns,
x"AA" after 21087000 ns,
x"E7" after 21098000 ns,
x"84" after 21109000 ns,
x"B7" after 21120000 ns,
x"17" after 21131000 ns,
x"00" after 21142000 ns,
x"00" after 21153000 ns,
x"83" after 21164000 ns,
x"A7" after 21175000 ns,
x"47" after 21186000 ns,
x"85" after 21197000 ns,
x"63" after 21208000 ns,
x"D8" after 21219000 ns,
x"07" after 21230000 ns,
x"00" after 21241000 ns,
x"B7" after 21252000 ns,
x"17" after 21263000 ns,
x"00" after 21274000 ns,
x"00" after 21285000 ns,
x"13" after 21296000 ns,
x"07" after 21307000 ns,
x"30" after 21318000 ns,
x"06" after 21329000 ns,
x"23" after 21340000 ns,
x"AA" after 21351000 ns,
x"E7" after 21362000 ns,
x"84" after 21373000 ns,
x"B7" after 21384000 ns,
x"17" after 21395000 ns,
x"00" after 21406000 ns,
x"00" after 21417000 ns,
x"03" after 21428000 ns,
x"A7" after 21439000 ns,
x"47" after 21450000 ns,
x"85" after 21461000 ns,
x"93" after 21472000 ns,
x"07" after 21483000 ns,
x"A0" after 21494000 ns,
x"00" after 21505000 ns,
x"33" after 21516000 ns,
x"47" after 21527000 ns,
x"F7" after 21538000 ns,
x"02" after 21549000 ns,
x"B7" after 21560000 ns,
x"17" after 21571000 ns,
x"00" after 21582000 ns,
x"00" after 21593000 ns,
x"93" after 21604000 ns,
x"87" after 21615000 ns,
x"07" after 21626000 ns,
x"80" after 21637000 ns,
x"23" after 21648000 ns,
x"A4" after 21659000 ns,
x"E7" after 21670000 ns,
x"00" after 21681000 ns,
x"B7" after 21692000 ns,
x"17" after 21703000 ns,
x"00" after 21714000 ns,
x"00" after 21725000 ns,
x"03" after 21736000 ns,
x"A7" after 21747000 ns,
x"47" after 21758000 ns,
x"85" after 21769000 ns,
x"93" after 21780000 ns,
x"07" after 21791000 ns,
x"A0" after 21802000 ns,
x"00" after 21813000 ns,
x"33" after 21824000 ns,
x"67" after 21835000 ns,
x"F7" after 21846000 ns,
x"02" after 21857000 ns,
x"B7" after 21868000 ns,
x"17" after 21879000 ns,
x"00" after 21890000 ns,
x"00" after 21901000 ns,
x"93" after 21912000 ns,
x"87" after 21923000 ns,
x"07" after 21934000 ns,
x"80" after 21945000 ns,
x"23" after 21956000 ns,
x"A6" after 21967000 ns,
x"E7" after 21978000 ns,
x"00" after 21989000 ns,
x"13" after 22000000 ns,
x"00" after 22011000 ns,
x"00" after 22022000 ns,
x"00" after 22033000 ns,
x"03" after 22044000 ns,
x"24" after 22055000 ns,
x"C1" after 22066000 ns,
x"00" after 22077000 ns,
x"13" after 22088000 ns,
x"01" after 22099000 ns,
x"01" after 22110000 ns,
x"01" after 22121000 ns,
x"67" after 22132000 ns,
x"80" after 22143000 ns,
x"00" after 22154000 ns,
x"00" after 22165000 ns,
x"13" after 22176000 ns,
x"01" after 22187000 ns,
x"01" after 22198000 ns,
x"FF" after 22209000 ns,
x"23" after 22220000 ns,
x"26" after 22231000 ns,
x"11" after 22242000 ns,
x"00" after 22253000 ns,
x"23" after 22264000 ns,
x"24" after 22275000 ns,
x"81" after 22286000 ns,
x"00" after 22297000 ns,
x"13" after 22308000 ns,
x"04" after 22319000 ns,
x"01" after 22330000 ns,
x"01" after 22341000 ns,
x"23" after 22352000 ns,
x"2A" after 22363000 ns,
x"04" after 22374000 ns,
x"FE" after 22385000 ns,
x"B7" after 22396000 ns,
x"17" after 22407000 ns,
x"00" after 22418000 ns,
x"00" after 22429000 ns,
x"13" after 22440000 ns,
x"85" after 22451000 ns,
x"C7" after 22462000 ns,
x"86" after 22473000 ns,
x"EF" after 22484000 ns,
x"F0" after 22495000 ns,
x"5F" after 22506000 ns,
x"8A" after 22517000 ns,
x"B7" after 22528000 ns,
x"67" after 22539000 ns,
x"00" after 22550000 ns,
x"80" after 22561000 ns,
x"37" after 22572000 ns,
x"C7" after 22583000 ns,
x"00" after 22594000 ns,
x"00" after 22605000 ns,
x"13" after 22616000 ns,
x"07" after 22627000 ns,
x"07" after 22638000 ns,
x"35" after 22649000 ns,
x"23" after 22660000 ns,
x"A0" after 22671000 ns,
x"E7" after 22682000 ns,
x"00" after 22693000 ns,
x"B7" after 22704000 ns,
x"67" after 22715000 ns,
x"00" after 22726000 ns,
x"80" after 22737000 ns,
x"93" after 22748000 ns,
x"87" after 22759000 ns,
x"07" after 22770000 ns,
x"01" after 22781000 ns,
x"13" after 22792000 ns,
x"07" after 22803000 ns,
x"A0" after 22814000 ns,
x"00" after 22825000 ns,
x"23" after 22836000 ns,
x"A0" after 22847000 ns,
x"E7" after 22858000 ns,
x"00" after 22869000 ns,
x"B7" after 22880000 ns,
x"67" after 22891000 ns,
x"00" after 22902000 ns,
x"80" after 22913000 ns,
x"93" after 22924000 ns,
x"87" after 22935000 ns,
x"07" after 22946000 ns,
x"02" after 22957000 ns,
x"13" after 22968000 ns,
x"07" after 22979000 ns,
x"10" after 22990000 ns,
x"00" after 23001000 ns,
x"23" after 23012000 ns,
x"80" after 23023000 ns,
x"E7" after 23034000 ns,
x"00" after 23045000 ns,
x"13" after 23056000 ns,
x"00" after 23067000 ns,
x"00" after 23078000 ns,
x"00" after 23089000 ns,
x"83" after 23100000 ns,
x"20" after 23111000 ns,
x"C1" after 23122000 ns,
x"00" after 23133000 ns,
x"03" after 23144000 ns,
x"24" after 23155000 ns,
x"81" after 23166000 ns,
x"00" after 23177000 ns,
x"13" after 23188000 ns,
x"01" after 23199000 ns,
x"01" after 23210000 ns,
x"01" after 23221000 ns,
x"67" after 23232000 ns,
x"80" after 23243000 ns,
x"00" after 23254000 ns,
x"00" after 23265000 ns,
x"13" after 23276000 ns,
x"01" after 23287000 ns,
x"01" after 23298000 ns,
x"FE" after 23309000 ns,
x"23" after 23320000 ns,
x"2E" after 23331000 ns,
x"11" after 23342000 ns,
x"00" after 23353000 ns,
x"23" after 23364000 ns,
x"2C" after 23375000 ns,
x"81" after 23386000 ns,
x"00" after 23397000 ns,
x"13" after 23408000 ns,
x"04" after 23419000 ns,
x"01" after 23430000 ns,
x"02" after 23441000 ns,
x"B7" after 23452000 ns,
x"07" after 23463000 ns,
x"00" after 23474000 ns,
x"FF" after 23485000 ns,
x"23" after 23496000 ns,
x"28" after 23507000 ns,
x"F4" after 23518000 ns,
x"FE" after 23529000 ns,
x"93" after 23540000 ns,
x"07" after 23551000 ns,
x"F0" after 23562000 ns,
x"FF" after 23573000 ns,
x"23" after 23584000 ns,
x"26" after 23595000 ns,
x"F4" after 23606000 ns,
x"FE" after 23617000 ns,
x"B7" after 23628000 ns,
x"07" after 23639000 ns,
x"00" after 23650000 ns,
x"C0" after 23661000 ns,
x"23" after 23672000 ns,
x"24" after 23683000 ns,
x"F4" after 23694000 ns,
x"FE" after 23705000 ns,
x"03" after 23716000 ns,
x"26" after 23727000 ns,
x"84" after 23738000 ns,
x"FE" after 23749000 ns,
x"83" after 23760000 ns,
x"25" after 23771000 ns,
x"C4" after 23782000 ns,
x"FE" after 23793000 ns,
x"03" after 23804000 ns,
x"25" after 23815000 ns,
x"04" after 23826000 ns,
x"FF" after 23837000 ns,
x"EF" after 23848000 ns,
x"F0" after 23859000 ns,
x"8F" after 23870000 ns,
x"FF" after 23881000 ns,
x"B7" after 23892000 ns,
x"17" after 23903000 ns,
x"00" after 23914000 ns,
x"00" after 23925000 ns,
x"13" after 23936000 ns,
x"85" after 23947000 ns,
x"87" after 23958000 ns,
x"87" after 23969000 ns,
x"EF" after 23980000 ns,
x"F0" after 23991000 ns,
x"DF" after 24002000 ns,
x"81" after 24013000 ns,
x"B7" after 24024000 ns,
x"27" after 24035000 ns,
x"00" after 24046000 ns,
x"00" after 24057000 ns,
x"93" after 24068000 ns,
x"85" after 24079000 ns,
x"C7" after 24090000 ns,
x"1D" after 24101000 ns,
x"13" after 24112000 ns,
x"05" after 24123000 ns,
x"10" after 24134000 ns,
x"00" after 24145000 ns,
x"EF" after 24156000 ns,
x"F0" after 24167000 ns,
x"CF" after 24178000 ns,
x"FA" after 24189000 ns,
x"B7" after 24200000 ns,
x"27" after 24211000 ns,
x"00" after 24222000 ns,
x"00" after 24233000 ns,
x"93" after 24244000 ns,
x"85" after 24255000 ns,
x"87" after 24266000 ns,
x"3A" after 24277000 ns,
x"13" after 24288000 ns,
x"05" after 24299000 ns,
x"70" after 24310000 ns,
x"00" after 24321000 ns,
x"EF" after 24332000 ns,
x"F0" after 24343000 ns,
x"CF" after 24354000 ns,
x"F9" after 24365000 ns,
x"B7" after 24376000 ns,
x"27" after 24387000 ns,
x"00" after 24398000 ns,
x"00" after 24409000 ns,
x"93" after 24420000 ns,
x"85" after 24431000 ns,
x"47" after 24442000 ns,
x"30" after 24453000 ns,
x"13" after 24464000 ns,
x"05" after 24475000 ns,
x"60" after 24486000 ns,
x"00" after 24497000 ns,
x"EF" after 24508000 ns,
x"F0" after 24519000 ns,
x"CF" after 24530000 ns,
x"F8" after 24541000 ns,
x"B7" after 24552000 ns,
x"17" after 24563000 ns,
x"00" after 24574000 ns,
x"00" after 24585000 ns,
x"13" after 24596000 ns,
x"85" after 24607000 ns,
x"87" after 24618000 ns,
x"88" after 24629000 ns,
x"EF" after 24640000 ns,
x"F0" after 24651000 ns,
x"0F" after 24662000 ns,
x"FE" after 24673000 ns,
x"13" after 24684000 ns,
x"05" after 24695000 ns,
x"30" after 24706000 ns,
x"0C" after 24717000 ns,
x"EF" after 24728000 ns,
x"F0" after 24739000 ns,
x"CF" after 24750000 ns,
x"FC" after 24761000 ns,
x"B7" after 24772000 ns,
x"17" after 24783000 ns,
x"00" after 24794000 ns,
x"00" after 24805000 ns,
x"13" after 24816000 ns,
x"85" after 24827000 ns,
x"07" after 24838000 ns,
x"8A" after 24849000 ns,
x"EF" after 24860000 ns,
x"F0" after 24871000 ns,
x"CF" after 24882000 ns,
x"FC" after 24893000 ns,
x"B7" after 24904000 ns,
x"C7" after 24915000 ns,
x"00" after 24926000 ns,
x"00" after 24937000 ns,
x"13" after 24948000 ns,
x"85" after 24959000 ns,
x"07" after 24970000 ns,
x"35" after 24981000 ns,
x"EF" after 24992000 ns,
x"F0" after 25003000 ns,
x"CF" after 25014000 ns,
x"F6" after 25025000 ns,
x"13" after 25036000 ns,
x"05" after 25047000 ns,
x"00" after 25058000 ns,
x"01" after 25069000 ns,
x"EF" after 25080000 ns,
x"F0" after 25091000 ns,
x"0F" after 25102000 ns,
x"F7" after 25113000 ns,
x"13" after 25124000 ns,
x"05" after 25135000 ns,
x"10" after 25146000 ns,
x"00" after 25157000 ns,
x"EF" after 25168000 ns,
x"F0" after 25179000 ns,
x"4F" after 25190000 ns,
x"F7" after 25201000 ns,
x"B7" after 25212000 ns,
x"17" after 25223000 ns,
x"00" after 25234000 ns,
x"00" after 25245000 ns,
x"13" after 25256000 ns,
x"85" after 25267000 ns,
x"C7" after 25278000 ns,
x"8A" after 25289000 ns,
x"EF" after 25300000 ns,
x"F0" after 25311000 ns,
x"4F" after 25322000 ns,
x"FA" after 25333000 ns,
x"23" after 25344000 ns,
x"2A" after 25355000 ns,
x"04" after 25366000 ns,
x"FE" after 25377000 ns,
x"23" after 25388000 ns,
x"22" after 25399000 ns,
x"04" after 25410000 ns,
x"FE" after 25421000 ns,
x"93" after 25432000 ns,
x"07" after 25443000 ns,
x"44" after 25454000 ns,
x"FE" after 25465000 ns,
x"13" after 25476000 ns,
x"85" after 25487000 ns,
x"07" after 25498000 ns,
x"00" after 25509000 ns,
x"EF" after 25520000 ns,
x"F0" after 25531000 ns,
x"8F" after 25542000 ns,
x"FA" after 25553000 ns,
x"93" after 25564000 ns,
x"07" after 25575000 ns,
x"05" after 25586000 ns,
x"00" after 25597000 ns,
x"63" after 25608000 ns,
x"88" after 25619000 ns,
x"07" after 25630000 ns,
x"00" after 25641000 ns,
x"83" after 25652000 ns,
x"27" after 25663000 ns,
x"44" after 25674000 ns,
x"FE" after 25685000 ns,
x"13" after 25696000 ns,
x"85" after 25707000 ns,
x"07" after 25718000 ns,
x"00" after 25729000 ns,
x"EF" after 25740000 ns,
x"F0" after 25751000 ns,
x"CF" after 25762000 ns,
x"F7" after 25773000 ns,
x"03" after 25784000 ns,
x"27" after 25795000 ns,
x"44" after 25806000 ns,
x"FF" after 25817000 ns,
x"B7" after 25828000 ns,
x"87" after 25839000 ns,
x"01" after 25850000 ns,
x"00" after 25861000 ns,
x"93" after 25872000 ns,
x"87" after 25883000 ns,
x"07" after 25894000 ns,
x"6A" after 25905000 ns,
x"63" after 25916000 ns,
x"D6" after 25927000 ns,
x"E7" after 25938000 ns,
x"06" after 25949000 ns,
x"23" after 25960000 ns,
x"2A" after 25971000 ns,
x"04" after 25982000 ns,
x"FE" after 25993000 ns,
x"B7" after 26004000 ns,
x"17" after 26015000 ns,
x"00" after 26026000 ns,
x"00" after 26037000 ns,
x"83" after 26048000 ns,
x"A7" after 26059000 ns,
x"07" after 26070000 ns,
x"85" after 26081000 ns,
x"13" after 26092000 ns,
x"87" after 26103000 ns,
x"17" after 26114000 ns,
x"00" after 26125000 ns,
x"B7" after 26136000 ns,
x"17" after 26147000 ns,
x"00" after 26158000 ns,
x"00" after 26169000 ns,
x"23" after 26180000 ns,
x"A8" after 26191000 ns,
x"E7" after 26202000 ns,
x"84" after 26213000 ns,
x"B7" after 26224000 ns,
x"17" after 26235000 ns,
x"00" after 26246000 ns,
x"00" after 26257000 ns,
x"03" after 26268000 ns,
x"A7" after 26279000 ns,
x"07" after 26290000 ns,
x"85" after 26301000 ns,
x"93" after 26312000 ns,
x"07" after 26323000 ns,
x"30" after 26334000 ns,
x"06" after 26345000 ns,
x"63" after 26356000 ns,
x"D6" after 26367000 ns,
x"E7" after 26378000 ns,
x"00" after 26389000 ns,
x"B7" after 26400000 ns,
x"17" after 26411000 ns,
x"00" after 26422000 ns,
x"00" after 26433000 ns,
x"23" after 26444000 ns,
x"A8" after 26455000 ns,
x"07" after 26466000 ns,
x"84" after 26477000 ns,
x"B7" after 26488000 ns,
x"17" after 26499000 ns,
x"00" after 26510000 ns,
x"00" after 26521000 ns,
x"03" after 26532000 ns,
x"A7" after 26543000 ns,
x"07" after 26554000 ns,
x"85" after 26565000 ns,
x"93" after 26576000 ns,
x"07" after 26587000 ns,
x"A0" after 26598000 ns,
x"00" after 26609000 ns,
x"33" after 26620000 ns,
x"47" after 26631000 ns,
x"F7" after 26642000 ns,
x"02" after 26653000 ns,
x"B7" after 26664000 ns,
x"17" after 26675000 ns,
x"00" after 26686000 ns,
x"00" after 26697000 ns,
x"93" after 26708000 ns,
x"87" after 26719000 ns,
x"07" after 26730000 ns,
x"80" after 26741000 ns,
x"23" after 26752000 ns,
x"A0" after 26763000 ns,
x"E7" after 26774000 ns,
x"00" after 26785000 ns,
x"B7" after 26796000 ns,
x"17" after 26807000 ns,
x"00" after 26818000 ns,
x"00" after 26829000 ns,
x"03" after 26840000 ns,
x"A7" after 26851000 ns,
x"07" after 26862000 ns,
x"85" after 26873000 ns,
x"93" after 26884000 ns,
x"07" after 26895000 ns,
x"A0" after 26906000 ns,
x"00" after 26917000 ns,
x"33" after 26928000 ns,
x"67" after 26939000 ns,
x"F7" after 26950000 ns,
x"02" after 26961000 ns,
x"B7" after 26972000 ns,
x"17" after 26983000 ns,
x"00" after 26994000 ns,
x"00" after 27005000 ns,
x"93" after 27016000 ns,
x"87" after 27027000 ns,
x"07" after 27038000 ns,
x"80" after 27049000 ns,
x"23" after 27060000 ns,
x"A2" after 27071000 ns,
x"E7" after 27082000 ns,
x"00" after 27093000 ns,
x"83" after 27104000 ns,
x"27" after 27115000 ns,
x"44" after 27126000 ns,
x"FF" after 27137000 ns,
x"93" after 27148000 ns,
x"87" after 27159000 ns,
x"17" after 27170000 ns,
x"00" after 27181000 ns,
x"23" after 27192000 ns,
x"2A" after 27203000 ns,
x"F4" after 27214000 ns,
x"FE" after 27225000 ns,
x"6F" after 27236000 ns,
x"F0" after 27247000 ns,
x"9F" after 27258000 ns,
x"F5" after 27269000 ns,
x"00" after 27280000 ns,
x"00" after 27291000 ns,
x"00" after 27302000 ns,
x"B9" after 27313000 ns,
x"00" after 27324000 ns,
x"00" after 27335000 ns,
x"00" after 27346000 ns,
x"00" after 27357000 ns,
x"00" after 27368000 ns,
x"00" after 27379000 ns,
x"00" after 27390000 ns,
x"00" after 27401000 ns,
x"00" after 27412000 ns,
x"00" after 27423000 ns,
x"00" after 27434000 ns,
x"00" after 27445000 ns,
x"00" after 27456000 ns,
x"00" after 27467000 ns,
x"00" after 27478000 ns,
x"00" after 27489000 ns,
x"00" after 27500000 ns,
x"0C" after 27511000 ns,
x"00" after 27522000 ns,
x"00" after 27533000 ns,
x"90" after 27544000 ns,
x"0F" after 27555000 ns,
x"00" after 27566000 ns,
x"00" after 27577000 ns,
x"40" after 27588000 ns,
x"0A" after 27599000 ns,
x"00" after 27610000 ns,
x"00" after 27621000 ns,
x"00" after 27632000 ns,
x"0B" after 27643000 ns,
x"00" after 27654000 ns,
x"00" after 27665000 ns,
x"90" after 27676000 ns,
x"09" after 27687000 ns,
x"00" after 27698000 ns,
x"00" after 27709000 ns,
x"20" after 27720000 ns,
x"09" after 27731000 ns,
x"00" after 27742000 ns,
x"00" after 27753000 ns,
x"20" after 27764000 ns,
x"08" after 27775000 ns,
x"00" after 27786000 ns,
x"00" after 27797000 ns,
x"80" after 27808000 ns,
x"0F" after 27819000 ns,
x"00" after 27830000 ns,
x"00" after 27841000 ns,
x"00" after 27852000 ns,
x"08" after 27863000 ns,
x"00" after 27874000 ns,
x"00" after 27885000 ns,
x"00" after 27896000 ns,
x"09" after 27907000 ns,
x"00" after 27918000 ns,
x"00" after 27929000 ns,
x"00" after 27940000 ns,
x"0A" after 27951000 ns,
x"00" after 27962000 ns,
x"00" after 27973000 ns,
x"30" after 27984000 ns,
x"08" after 27995000 ns,
x"00" after 28006000 ns,
x"00" after 28017000 ns,
x"60" after 28028000 ns,
x"0C" after 28039000 ns,
x"00" after 28050000 ns,
x"00" after 28061000 ns,
x"10" after 28072000 ns,
x"0A" after 28083000 ns,
x"00" after 28094000 ns,
x"00" after 28105000 ns,
x"60" after 28116000 ns,
x"08" after 28127000 ns,
x"00" after 28138000 ns,
x"00" after 28149000 ns,
x"E0" after 28160000 ns,
x"08" after 28171000 ns,
x"00" after 28182000 ns,
x"00" after 28193000 ns,
x"00" after 28204000 ns,
x"00" after 28215000 ns,
x"00" after 28226000 ns,
x"00" after 28237000 ns,
x"00" after 28248000 ns,
x"00" after 28259000 ns,
x"00" after 28270000 ns,
x"00" after 28281000 ns,
x"30" after 28292000 ns,
x"31" after 28303000 ns,
x"32" after 28314000 ns,
x"33" after 28325000 ns,
x"34" after 28336000 ns,
x"35" after 28347000 ns,
x"36" after 28358000 ns,
x"37" after 28369000 ns,
x"38" after 28380000 ns,
x"39" after 28391000 ns,
x"41" after 28402000 ns,
x"42" after 28413000 ns,
x"43" after 28424000 ns,
x"44" after 28435000 ns,
x"45" after 28446000 ns,
x"46" after 28457000 ns,
x"00" after 28468000 ns,
x"00" after 28479000 ns,
x"00" after 28490000 ns,
x"00" after 28501000 ns,
x"43" after 28512000 ns,
x"61" after 28523000 ns,
x"6C" after 28534000 ns,
x"6C" after 28545000 ns,
x"5F" after 28556000 ns,
x"44" after 28567000 ns,
x"39" after 28578000 ns,
x"0A" after 28589000 ns,
x"00" after 28600000 ns,
x"00" after 28611000 ns,
x"00" after 28622000 ns,
x"00" after 28633000 ns,
x"53" after 28644000 ns,
x"45" after 28655000 ns,
x"54" after 28666000 ns,
x"55" after 28677000 ns,
x"50" after 28688000 ns,
x"20" after 28699000 ns,
x"42" after 28710000 ns,
x"44" after 28721000 ns,
x"20" after 28732000 ns,
x"50" after 28743000 ns,
x"4F" after 28754000 ns,
x"52" after 28765000 ns,
x"54" after 28776000 ns,
x"0A" after 28787000 ns,
x"00" after 28798000 ns,
x"00" after 28809000 ns,
x"53" after 28820000 ns,
x"45" after 28831000 ns,
x"54" after 28842000 ns,
x"55" after 28853000 ns,
x"50" after 28864000 ns,
x"20" after 28875000 ns,
x"54" after 28886000 ns,
x"49" after 28897000 ns,
x"4D" after 28908000 ns,
x"45" after 28919000 ns,
x"52" after 28930000 ns,
x"20" after 28941000 ns,
x"43" after 28952000 ns,
x"41" after 28963000 ns,
x"4C" after 28974000 ns,
x"4C" after 28985000 ns,
x"42" after 28996000 ns,
x"41" after 29007000 ns,
x"43" after 29018000 ns,
x"4B" after 29029000 ns,
x"20" after 29040000 ns,
x"0A" after 29051000 ns,
x"00" after 29062000 ns,
x"00" after 29073000 ns,
x"53" after 29084000 ns,
x"45" after 29095000 ns,
x"54" after 29106000 ns,
x"55" after 29117000 ns,
x"50" after 29128000 ns,
x"20" after 29139000 ns,
x"50" after 29150000 ns,
x"49" after 29161000 ns,
x"43" after 29172000 ns,
x"20" after 29183000 ns,
x"0A" after 29194000 ns,
x"00" after 29205000 ns,
x"53" after 29216000 ns,
x"45" after 29227000 ns,
x"54" after 29238000 ns,
x"55" after 29249000 ns,
x"50" after 29260000 ns,
x"20" after 29271000 ns,
x"54" after 29282000 ns,
x"49" after 29293000 ns,
x"4D" after 29304000 ns,
x"45" after 29315000 ns,
x"52" after 29326000 ns,
x"0A" after 29337000 ns,
x"00" after 29348000 ns;

-- VHDL for tx_dv:
tx_dv <= '1' after 0 ns, '0' after 50 ns,
'1' after 11000 ns, '0' after 11050 ns,
'1' after 22000 ns, '0' after 22050 ns,
'1' after 33000 ns, '0' after 33050 ns,
'1' after 44000 ns, '0' after 44050 ns,
'1' after 55000 ns, '0' after 55050 ns,
'1' after 66000 ns, '0' after 66050 ns,
'1' after 77000 ns, '0' after 77050 ns,
'1' after 88000 ns, '0' after 88050 ns,
'1' after 99000 ns, '0' after 99050 ns,
'1' after 110000 ns, '0' after 110050 ns,
'1' after 121000 ns, '0' after 121050 ns,
'1' after 132000 ns, '0' after 132050 ns,
'1' after 143000 ns, '0' after 143050 ns,
'1' after 154000 ns, '0' after 154050 ns,
'1' after 165000 ns, '0' after 165050 ns,
'1' after 176000 ns, '0' after 176050 ns,
'1' after 187000 ns, '0' after 187050 ns,
'1' after 198000 ns, '0' after 198050 ns,
'1' after 209000 ns, '0' after 209050 ns,
'1' after 220000 ns, '0' after 220050 ns,
'1' after 231000 ns, '0' after 231050 ns,
'1' after 242000 ns, '0' after 242050 ns,
'1' after 253000 ns, '0' after 253050 ns,
'1' after 264000 ns, '0' after 264050 ns,
'1' after 275000 ns, '0' after 275050 ns,
'1' after 286000 ns, '0' after 286050 ns,
'1' after 297000 ns, '0' after 297050 ns,
'1' after 308000 ns, '0' after 308050 ns,
'1' after 319000 ns, '0' after 319050 ns,
'1' after 330000 ns, '0' after 330050 ns,
'1' after 341000 ns, '0' after 341050 ns,
'1' after 352000 ns, '0' after 352050 ns,
'1' after 363000 ns, '0' after 363050 ns,
'1' after 374000 ns, '0' after 374050 ns,
'1' after 385000 ns, '0' after 385050 ns,
'1' after 396000 ns, '0' after 396050 ns,
'1' after 407000 ns, '0' after 407050 ns,
'1' after 418000 ns, '0' after 418050 ns,
'1' after 429000 ns, '0' after 429050 ns,
'1' after 440000 ns, '0' after 440050 ns,
'1' after 451000 ns, '0' after 451050 ns,
'1' after 462000 ns, '0' after 462050 ns,
'1' after 473000 ns, '0' after 473050 ns,
'1' after 484000 ns, '0' after 484050 ns,
'1' after 495000 ns, '0' after 495050 ns,
'1' after 506000 ns, '0' after 506050 ns,
'1' after 517000 ns, '0' after 517050 ns,
'1' after 528000 ns, '0' after 528050 ns,
'1' after 539000 ns, '0' after 539050 ns,
'1' after 550000 ns, '0' after 550050 ns,
'1' after 561000 ns, '0' after 561050 ns,
'1' after 572000 ns, '0' after 572050 ns,
'1' after 583000 ns, '0' after 583050 ns,
'1' after 594000 ns, '0' after 594050 ns,
'1' after 605000 ns, '0' after 605050 ns,
'1' after 616000 ns, '0' after 616050 ns,
'1' after 627000 ns, '0' after 627050 ns,
'1' after 638000 ns, '0' after 638050 ns,
'1' after 649000 ns, '0' after 649050 ns,
'1' after 660000 ns, '0' after 660050 ns,
'1' after 671000 ns, '0' after 671050 ns,
'1' after 682000 ns, '0' after 682050 ns,
'1' after 693000 ns, '0' after 693050 ns,
'1' after 704000 ns, '0' after 704050 ns,
'1' after 715000 ns, '0' after 715050 ns,
'1' after 726000 ns, '0' after 726050 ns,
'1' after 737000 ns, '0' after 737050 ns,
'1' after 748000 ns, '0' after 748050 ns,
'1' after 759000 ns, '0' after 759050 ns,
'1' after 770000 ns, '0' after 770050 ns,
'1' after 781000 ns, '0' after 781050 ns,
'1' after 792000 ns, '0' after 792050 ns,
'1' after 803000 ns, '0' after 803050 ns,
'1' after 814000 ns, '0' after 814050 ns,
'1' after 825000 ns, '0' after 825050 ns,
'1' after 836000 ns, '0' after 836050 ns,
'1' after 847000 ns, '0' after 847050 ns,
'1' after 858000 ns, '0' after 858050 ns,
'1' after 869000 ns, '0' after 869050 ns,
'1' after 880000 ns, '0' after 880050 ns,
'1' after 891000 ns, '0' after 891050 ns,
'1' after 902000 ns, '0' after 902050 ns,
'1' after 913000 ns, '0' after 913050 ns,
'1' after 924000 ns, '0' after 924050 ns,
'1' after 935000 ns, '0' after 935050 ns,
'1' after 946000 ns, '0' after 946050 ns,
'1' after 957000 ns, '0' after 957050 ns,
'1' after 968000 ns, '0' after 968050 ns,
'1' after 979000 ns, '0' after 979050 ns,
'1' after 990000 ns, '0' after 990050 ns,
'1' after 1001000 ns, '0' after 1001050 ns,
'1' after 1012000 ns, '0' after 1012050 ns,
'1' after 1023000 ns, '0' after 1023050 ns,
'1' after 1034000 ns, '0' after 1034050 ns,
'1' after 1045000 ns, '0' after 1045050 ns,
'1' after 1056000 ns, '0' after 1056050 ns,
'1' after 1067000 ns, '0' after 1067050 ns,
'1' after 1078000 ns, '0' after 1078050 ns,
'1' after 1089000 ns, '0' after 1089050 ns,
'1' after 1100000 ns, '0' after 1100050 ns,
'1' after 1111000 ns, '0' after 1111050 ns,
'1' after 1122000 ns, '0' after 1122050 ns,
'1' after 1133000 ns, '0' after 1133050 ns,
'1' after 1144000 ns, '0' after 1144050 ns,
'1' after 1155000 ns, '0' after 1155050 ns,
'1' after 1166000 ns, '0' after 1166050 ns,
'1' after 1177000 ns, '0' after 1177050 ns,
'1' after 1188000 ns, '0' after 1188050 ns,
'1' after 1199000 ns, '0' after 1199050 ns,
'1' after 1210000 ns, '0' after 1210050 ns,
'1' after 1221000 ns, '0' after 1221050 ns,
'1' after 1232000 ns, '0' after 1232050 ns,
'1' after 1243000 ns, '0' after 1243050 ns,
'1' after 1254000 ns, '0' after 1254050 ns,
'1' after 1265000 ns, '0' after 1265050 ns,
'1' after 1276000 ns, '0' after 1276050 ns,
'1' after 1287000 ns, '0' after 1287050 ns,
'1' after 1298000 ns, '0' after 1298050 ns,
'1' after 1309000 ns, '0' after 1309050 ns,
'1' after 1320000 ns, '0' after 1320050 ns,
'1' after 1331000 ns, '0' after 1331050 ns,
'1' after 1342000 ns, '0' after 1342050 ns,
'1' after 1353000 ns, '0' after 1353050 ns,
'1' after 1364000 ns, '0' after 1364050 ns,
'1' after 1375000 ns, '0' after 1375050 ns,
'1' after 1386000 ns, '0' after 1386050 ns,
'1' after 1397000 ns, '0' after 1397050 ns,
'1' after 1408000 ns, '0' after 1408050 ns,
'1' after 1419000 ns, '0' after 1419050 ns,
'1' after 1430000 ns, '0' after 1430050 ns,
'1' after 1441000 ns, '0' after 1441050 ns,
'1' after 1452000 ns, '0' after 1452050 ns,
'1' after 1463000 ns, '0' after 1463050 ns,
'1' after 1474000 ns, '0' after 1474050 ns,
'1' after 1485000 ns, '0' after 1485050 ns,
'1' after 1496000 ns, '0' after 1496050 ns,
'1' after 1507000 ns, '0' after 1507050 ns,
'1' after 1518000 ns, '0' after 1518050 ns,
'1' after 1529000 ns, '0' after 1529050 ns,
'1' after 1540000 ns, '0' after 1540050 ns,
'1' after 1551000 ns, '0' after 1551050 ns,
'1' after 1562000 ns, '0' after 1562050 ns,
'1' after 1573000 ns, '0' after 1573050 ns,
'1' after 1584000 ns, '0' after 1584050 ns,
'1' after 1595000 ns, '0' after 1595050 ns,
'1' after 1606000 ns, '0' after 1606050 ns,
'1' after 1617000 ns, '0' after 1617050 ns,
'1' after 1628000 ns, '0' after 1628050 ns,
'1' after 1639000 ns, '0' after 1639050 ns,
'1' after 1650000 ns, '0' after 1650050 ns,
'1' after 1661000 ns, '0' after 1661050 ns,
'1' after 1672000 ns, '0' after 1672050 ns,
'1' after 1683000 ns, '0' after 1683050 ns,
'1' after 1694000 ns, '0' after 1694050 ns,
'1' after 1705000 ns, '0' after 1705050 ns,
'1' after 1716000 ns, '0' after 1716050 ns,
'1' after 1727000 ns, '0' after 1727050 ns,
'1' after 1738000 ns, '0' after 1738050 ns,
'1' after 1749000 ns, '0' after 1749050 ns,
'1' after 1760000 ns, '0' after 1760050 ns,
'1' after 1771000 ns, '0' after 1771050 ns,
'1' after 1782000 ns, '0' after 1782050 ns,
'1' after 1793000 ns, '0' after 1793050 ns,
'1' after 1804000 ns, '0' after 1804050 ns,
'1' after 1815000 ns, '0' after 1815050 ns,
'1' after 1826000 ns, '0' after 1826050 ns,
'1' after 1837000 ns, '0' after 1837050 ns,
'1' after 1848000 ns, '0' after 1848050 ns,
'1' after 1859000 ns, '0' after 1859050 ns,
'1' after 1870000 ns, '0' after 1870050 ns,
'1' after 1881000 ns, '0' after 1881050 ns,
'1' after 1892000 ns, '0' after 1892050 ns,
'1' after 1903000 ns, '0' after 1903050 ns,
'1' after 1914000 ns, '0' after 1914050 ns,
'1' after 1925000 ns, '0' after 1925050 ns,
'1' after 1936000 ns, '0' after 1936050 ns,
'1' after 1947000 ns, '0' after 1947050 ns,
'1' after 1958000 ns, '0' after 1958050 ns,
'1' after 1969000 ns, '0' after 1969050 ns,
'1' after 1980000 ns, '0' after 1980050 ns,
'1' after 1991000 ns, '0' after 1991050 ns,
'1' after 2002000 ns, '0' after 2002050 ns,
'1' after 2013000 ns, '0' after 2013050 ns,
'1' after 2024000 ns, '0' after 2024050 ns,
'1' after 2035000 ns, '0' after 2035050 ns,
'1' after 2046000 ns, '0' after 2046050 ns,
'1' after 2057000 ns, '0' after 2057050 ns,
'1' after 2068000 ns, '0' after 2068050 ns,
'1' after 2079000 ns, '0' after 2079050 ns,
'1' after 2090000 ns, '0' after 2090050 ns,
'1' after 2101000 ns, '0' after 2101050 ns,
'1' after 2112000 ns, '0' after 2112050 ns,
'1' after 2123000 ns, '0' after 2123050 ns,
'1' after 2134000 ns, '0' after 2134050 ns,
'1' after 2145000 ns, '0' after 2145050 ns,
'1' after 2156000 ns, '0' after 2156050 ns,
'1' after 2167000 ns, '0' after 2167050 ns,
'1' after 2178000 ns, '0' after 2178050 ns,
'1' after 2189000 ns, '0' after 2189050 ns,
'1' after 2200000 ns, '0' after 2200050 ns,
'1' after 2211000 ns, '0' after 2211050 ns,
'1' after 2222000 ns, '0' after 2222050 ns,
'1' after 2233000 ns, '0' after 2233050 ns,
'1' after 2244000 ns, '0' after 2244050 ns,
'1' after 2255000 ns, '0' after 2255050 ns,
'1' after 2266000 ns, '0' after 2266050 ns,
'1' after 2277000 ns, '0' after 2277050 ns,
'1' after 2288000 ns, '0' after 2288050 ns,
'1' after 2299000 ns, '0' after 2299050 ns,
'1' after 2310000 ns, '0' after 2310050 ns,
'1' after 2321000 ns, '0' after 2321050 ns,
'1' after 2332000 ns, '0' after 2332050 ns,
'1' after 2343000 ns, '0' after 2343050 ns,
'1' after 2354000 ns, '0' after 2354050 ns,
'1' after 2365000 ns, '0' after 2365050 ns,
'1' after 2376000 ns, '0' after 2376050 ns,
'1' after 2387000 ns, '0' after 2387050 ns,
'1' after 2398000 ns, '0' after 2398050 ns,
'1' after 2409000 ns, '0' after 2409050 ns,
'1' after 2420000 ns, '0' after 2420050 ns,
'1' after 2431000 ns, '0' after 2431050 ns,
'1' after 2442000 ns, '0' after 2442050 ns,
'1' after 2453000 ns, '0' after 2453050 ns,
'1' after 2464000 ns, '0' after 2464050 ns,
'1' after 2475000 ns, '0' after 2475050 ns,
'1' after 2486000 ns, '0' after 2486050 ns,
'1' after 2497000 ns, '0' after 2497050 ns,
'1' after 2508000 ns, '0' after 2508050 ns,
'1' after 2519000 ns, '0' after 2519050 ns,
'1' after 2530000 ns, '0' after 2530050 ns,
'1' after 2541000 ns, '0' after 2541050 ns,
'1' after 2552000 ns, '0' after 2552050 ns,
'1' after 2563000 ns, '0' after 2563050 ns,
'1' after 2574000 ns, '0' after 2574050 ns,
'1' after 2585000 ns, '0' after 2585050 ns,
'1' after 2596000 ns, '0' after 2596050 ns,
'1' after 2607000 ns, '0' after 2607050 ns,
'1' after 2618000 ns, '0' after 2618050 ns,
'1' after 2629000 ns, '0' after 2629050 ns,
'1' after 2640000 ns, '0' after 2640050 ns,
'1' after 2651000 ns, '0' after 2651050 ns,
'1' after 2662000 ns, '0' after 2662050 ns,
'1' after 2673000 ns, '0' after 2673050 ns,
'1' after 2684000 ns, '0' after 2684050 ns,
'1' after 2695000 ns, '0' after 2695050 ns,
'1' after 2706000 ns, '0' after 2706050 ns,
'1' after 2717000 ns, '0' after 2717050 ns,
'1' after 2728000 ns, '0' after 2728050 ns,
'1' after 2739000 ns, '0' after 2739050 ns,
'1' after 2750000 ns, '0' after 2750050 ns,
'1' after 2761000 ns, '0' after 2761050 ns,
'1' after 2772000 ns, '0' after 2772050 ns,
'1' after 2783000 ns, '0' after 2783050 ns,
'1' after 2794000 ns, '0' after 2794050 ns,
'1' after 2805000 ns, '0' after 2805050 ns,
'1' after 2816000 ns, '0' after 2816050 ns,
'1' after 2827000 ns, '0' after 2827050 ns,
'1' after 2838000 ns, '0' after 2838050 ns,
'1' after 2849000 ns, '0' after 2849050 ns,
'1' after 2860000 ns, '0' after 2860050 ns,
'1' after 2871000 ns, '0' after 2871050 ns,
'1' after 2882000 ns, '0' after 2882050 ns,
'1' after 2893000 ns, '0' after 2893050 ns,
'1' after 2904000 ns, '0' after 2904050 ns,
'1' after 2915000 ns, '0' after 2915050 ns,
'1' after 2926000 ns, '0' after 2926050 ns,
'1' after 2937000 ns, '0' after 2937050 ns,
'1' after 2948000 ns, '0' after 2948050 ns,
'1' after 2959000 ns, '0' after 2959050 ns,
'1' after 2970000 ns, '0' after 2970050 ns,
'1' after 2981000 ns, '0' after 2981050 ns,
'1' after 2992000 ns, '0' after 2992050 ns,
'1' after 3003000 ns, '0' after 3003050 ns,
'1' after 3014000 ns, '0' after 3014050 ns,
'1' after 3025000 ns, '0' after 3025050 ns,
'1' after 3036000 ns, '0' after 3036050 ns,
'1' after 3047000 ns, '0' after 3047050 ns,
'1' after 3058000 ns, '0' after 3058050 ns,
'1' after 3069000 ns, '0' after 3069050 ns,
'1' after 3080000 ns, '0' after 3080050 ns,
'1' after 3091000 ns, '0' after 3091050 ns,
'1' after 3102000 ns, '0' after 3102050 ns,
'1' after 3113000 ns, '0' after 3113050 ns,
'1' after 3124000 ns, '0' after 3124050 ns,
'1' after 3135000 ns, '0' after 3135050 ns,
'1' after 3146000 ns, '0' after 3146050 ns,
'1' after 3157000 ns, '0' after 3157050 ns,
'1' after 3168000 ns, '0' after 3168050 ns,
'1' after 3179000 ns, '0' after 3179050 ns,
'1' after 3190000 ns, '0' after 3190050 ns,
'1' after 3201000 ns, '0' after 3201050 ns,
'1' after 3212000 ns, '0' after 3212050 ns,
'1' after 3223000 ns, '0' after 3223050 ns,
'1' after 3234000 ns, '0' after 3234050 ns,
'1' after 3245000 ns, '0' after 3245050 ns,
'1' after 3256000 ns, '0' after 3256050 ns,
'1' after 3267000 ns, '0' after 3267050 ns,
'1' after 3278000 ns, '0' after 3278050 ns,
'1' after 3289000 ns, '0' after 3289050 ns,
'1' after 3300000 ns, '0' after 3300050 ns,
'1' after 3311000 ns, '0' after 3311050 ns,
'1' after 3322000 ns, '0' after 3322050 ns,
'1' after 3333000 ns, '0' after 3333050 ns,
'1' after 3344000 ns, '0' after 3344050 ns,
'1' after 3355000 ns, '0' after 3355050 ns,
'1' after 3366000 ns, '0' after 3366050 ns,
'1' after 3377000 ns, '0' after 3377050 ns,
'1' after 3388000 ns, '0' after 3388050 ns,
'1' after 3399000 ns, '0' after 3399050 ns,
'1' after 3410000 ns, '0' after 3410050 ns,
'1' after 3421000 ns, '0' after 3421050 ns,
'1' after 3432000 ns, '0' after 3432050 ns,
'1' after 3443000 ns, '0' after 3443050 ns,
'1' after 3454000 ns, '0' after 3454050 ns,
'1' after 3465000 ns, '0' after 3465050 ns,
'1' after 3476000 ns, '0' after 3476050 ns,
'1' after 3487000 ns, '0' after 3487050 ns,
'1' after 3498000 ns, '0' after 3498050 ns,
'1' after 3509000 ns, '0' after 3509050 ns,
'1' after 3520000 ns, '0' after 3520050 ns,
'1' after 3531000 ns, '0' after 3531050 ns,
'1' after 3542000 ns, '0' after 3542050 ns,
'1' after 3553000 ns, '0' after 3553050 ns,
'1' after 3564000 ns, '0' after 3564050 ns,
'1' after 3575000 ns, '0' after 3575050 ns,
'1' after 3586000 ns, '0' after 3586050 ns,
'1' after 3597000 ns, '0' after 3597050 ns,
'1' after 3608000 ns, '0' after 3608050 ns,
'1' after 3619000 ns, '0' after 3619050 ns,
'1' after 3630000 ns, '0' after 3630050 ns,
'1' after 3641000 ns, '0' after 3641050 ns,
'1' after 3652000 ns, '0' after 3652050 ns,
'1' after 3663000 ns, '0' after 3663050 ns,
'1' after 3674000 ns, '0' after 3674050 ns,
'1' after 3685000 ns, '0' after 3685050 ns,
'1' after 3696000 ns, '0' after 3696050 ns,
'1' after 3707000 ns, '0' after 3707050 ns,
'1' after 3718000 ns, '0' after 3718050 ns,
'1' after 3729000 ns, '0' after 3729050 ns,
'1' after 3740000 ns, '0' after 3740050 ns,
'1' after 3751000 ns, '0' after 3751050 ns,
'1' after 3762000 ns, '0' after 3762050 ns,
'1' after 3773000 ns, '0' after 3773050 ns,
'1' after 3784000 ns, '0' after 3784050 ns,
'1' after 3795000 ns, '0' after 3795050 ns,
'1' after 3806000 ns, '0' after 3806050 ns,
'1' after 3817000 ns, '0' after 3817050 ns,
'1' after 3828000 ns, '0' after 3828050 ns,
'1' after 3839000 ns, '0' after 3839050 ns,
'1' after 3850000 ns, '0' after 3850050 ns,
'1' after 3861000 ns, '0' after 3861050 ns,
'1' after 3872000 ns, '0' after 3872050 ns,
'1' after 3883000 ns, '0' after 3883050 ns,
'1' after 3894000 ns, '0' after 3894050 ns,
'1' after 3905000 ns, '0' after 3905050 ns,
'1' after 3916000 ns, '0' after 3916050 ns,
'1' after 3927000 ns, '0' after 3927050 ns,
'1' after 3938000 ns, '0' after 3938050 ns,
'1' after 3949000 ns, '0' after 3949050 ns,
'1' after 3960000 ns, '0' after 3960050 ns,
'1' after 3971000 ns, '0' after 3971050 ns,
'1' after 3982000 ns, '0' after 3982050 ns,
'1' after 3993000 ns, '0' after 3993050 ns,
'1' after 4004000 ns, '0' after 4004050 ns,
'1' after 4015000 ns, '0' after 4015050 ns,
'1' after 4026000 ns, '0' after 4026050 ns,
'1' after 4037000 ns, '0' after 4037050 ns,
'1' after 4048000 ns, '0' after 4048050 ns,
'1' after 4059000 ns, '0' after 4059050 ns,
'1' after 4070000 ns, '0' after 4070050 ns,
'1' after 4081000 ns, '0' after 4081050 ns,
'1' after 4092000 ns, '0' after 4092050 ns,
'1' after 4103000 ns, '0' after 4103050 ns,
'1' after 4114000 ns, '0' after 4114050 ns,
'1' after 4125000 ns, '0' after 4125050 ns,
'1' after 4136000 ns, '0' after 4136050 ns,
'1' after 4147000 ns, '0' after 4147050 ns,
'1' after 4158000 ns, '0' after 4158050 ns,
'1' after 4169000 ns, '0' after 4169050 ns,
'1' after 4180000 ns, '0' after 4180050 ns,
'1' after 4191000 ns, '0' after 4191050 ns,
'1' after 4202000 ns, '0' after 4202050 ns,
'1' after 4213000 ns, '0' after 4213050 ns,
'1' after 4224000 ns, '0' after 4224050 ns,
'1' after 4235000 ns, '0' after 4235050 ns,
'1' after 4246000 ns, '0' after 4246050 ns,
'1' after 4257000 ns, '0' after 4257050 ns,
'1' after 4268000 ns, '0' after 4268050 ns,
'1' after 4279000 ns, '0' after 4279050 ns,
'1' after 4290000 ns, '0' after 4290050 ns,
'1' after 4301000 ns, '0' after 4301050 ns,
'1' after 4312000 ns, '0' after 4312050 ns,
'1' after 4323000 ns, '0' after 4323050 ns,
'1' after 4334000 ns, '0' after 4334050 ns,
'1' after 4345000 ns, '0' after 4345050 ns,
'1' after 4356000 ns, '0' after 4356050 ns,
'1' after 4367000 ns, '0' after 4367050 ns,
'1' after 4378000 ns, '0' after 4378050 ns,
'1' after 4389000 ns, '0' after 4389050 ns,
'1' after 4400000 ns, '0' after 4400050 ns,
'1' after 4411000 ns, '0' after 4411050 ns,
'1' after 4422000 ns, '0' after 4422050 ns,
'1' after 4433000 ns, '0' after 4433050 ns,
'1' after 4444000 ns, '0' after 4444050 ns,
'1' after 4455000 ns, '0' after 4455050 ns,
'1' after 4466000 ns, '0' after 4466050 ns,
'1' after 4477000 ns, '0' after 4477050 ns,
'1' after 4488000 ns, '0' after 4488050 ns,
'1' after 4499000 ns, '0' after 4499050 ns,
'1' after 4510000 ns, '0' after 4510050 ns,
'1' after 4521000 ns, '0' after 4521050 ns,
'1' after 4532000 ns, '0' after 4532050 ns,
'1' after 4543000 ns, '0' after 4543050 ns,
'1' after 4554000 ns, '0' after 4554050 ns,
'1' after 4565000 ns, '0' after 4565050 ns,
'1' after 4576000 ns, '0' after 4576050 ns,
'1' after 4587000 ns, '0' after 4587050 ns,
'1' after 4598000 ns, '0' after 4598050 ns,
'1' after 4609000 ns, '0' after 4609050 ns,
'1' after 4620000 ns, '0' after 4620050 ns,
'1' after 4631000 ns, '0' after 4631050 ns,
'1' after 4642000 ns, '0' after 4642050 ns,
'1' after 4653000 ns, '0' after 4653050 ns,
'1' after 4664000 ns, '0' after 4664050 ns,
'1' after 4675000 ns, '0' after 4675050 ns,
'1' after 4686000 ns, '0' after 4686050 ns,
'1' after 4697000 ns, '0' after 4697050 ns,
'1' after 4708000 ns, '0' after 4708050 ns,
'1' after 4719000 ns, '0' after 4719050 ns,
'1' after 4730000 ns, '0' after 4730050 ns,
'1' after 4741000 ns, '0' after 4741050 ns,
'1' after 4752000 ns, '0' after 4752050 ns,
'1' after 4763000 ns, '0' after 4763050 ns,
'1' after 4774000 ns, '0' after 4774050 ns,
'1' after 4785000 ns, '0' after 4785050 ns,
'1' after 4796000 ns, '0' after 4796050 ns,
'1' after 4807000 ns, '0' after 4807050 ns,
'1' after 4818000 ns, '0' after 4818050 ns,
'1' after 4829000 ns, '0' after 4829050 ns,
'1' after 4840000 ns, '0' after 4840050 ns,
'1' after 4851000 ns, '0' after 4851050 ns,
'1' after 4862000 ns, '0' after 4862050 ns,
'1' after 4873000 ns, '0' after 4873050 ns,
'1' after 4884000 ns, '0' after 4884050 ns,
'1' after 4895000 ns, '0' after 4895050 ns,
'1' after 4906000 ns, '0' after 4906050 ns,
'1' after 4917000 ns, '0' after 4917050 ns,
'1' after 4928000 ns, '0' after 4928050 ns,
'1' after 4939000 ns, '0' after 4939050 ns,
'1' after 4950000 ns, '0' after 4950050 ns,
'1' after 4961000 ns, '0' after 4961050 ns,
'1' after 4972000 ns, '0' after 4972050 ns,
'1' after 4983000 ns, '0' after 4983050 ns,
'1' after 4994000 ns, '0' after 4994050 ns,
'1' after 5005000 ns, '0' after 5005050 ns,
'1' after 5016000 ns, '0' after 5016050 ns,
'1' after 5027000 ns, '0' after 5027050 ns,
'1' after 5038000 ns, '0' after 5038050 ns,
'1' after 5049000 ns, '0' after 5049050 ns,
'1' after 5060000 ns, '0' after 5060050 ns,
'1' after 5071000 ns, '0' after 5071050 ns,
'1' after 5082000 ns, '0' after 5082050 ns,
'1' after 5093000 ns, '0' after 5093050 ns,
'1' after 5104000 ns, '0' after 5104050 ns,
'1' after 5115000 ns, '0' after 5115050 ns,
'1' after 5126000 ns, '0' after 5126050 ns,
'1' after 5137000 ns, '0' after 5137050 ns,
'1' after 5148000 ns, '0' after 5148050 ns,
'1' after 5159000 ns, '0' after 5159050 ns,
'1' after 5170000 ns, '0' after 5170050 ns,
'1' after 5181000 ns, '0' after 5181050 ns,
'1' after 5192000 ns, '0' after 5192050 ns,
'1' after 5203000 ns, '0' after 5203050 ns,
'1' after 5214000 ns, '0' after 5214050 ns,
'1' after 5225000 ns, '0' after 5225050 ns,
'1' after 5236000 ns, '0' after 5236050 ns,
'1' after 5247000 ns, '0' after 5247050 ns,
'1' after 5258000 ns, '0' after 5258050 ns,
'1' after 5269000 ns, '0' after 5269050 ns,
'1' after 5280000 ns, '0' after 5280050 ns,
'1' after 5291000 ns, '0' after 5291050 ns,
'1' after 5302000 ns, '0' after 5302050 ns,
'1' after 5313000 ns, '0' after 5313050 ns,
'1' after 5324000 ns, '0' after 5324050 ns,
'1' after 5335000 ns, '0' after 5335050 ns,
'1' after 5346000 ns, '0' after 5346050 ns,
'1' after 5357000 ns, '0' after 5357050 ns,
'1' after 5368000 ns, '0' after 5368050 ns,
'1' after 5379000 ns, '0' after 5379050 ns,
'1' after 5390000 ns, '0' after 5390050 ns,
'1' after 5401000 ns, '0' after 5401050 ns,
'1' after 5412000 ns, '0' after 5412050 ns,
'1' after 5423000 ns, '0' after 5423050 ns,
'1' after 5434000 ns, '0' after 5434050 ns,
'1' after 5445000 ns, '0' after 5445050 ns,
'1' after 5456000 ns, '0' after 5456050 ns,
'1' after 5467000 ns, '0' after 5467050 ns,
'1' after 5478000 ns, '0' after 5478050 ns,
'1' after 5489000 ns, '0' after 5489050 ns,
'1' after 5500000 ns, '0' after 5500050 ns,
'1' after 5511000 ns, '0' after 5511050 ns,
'1' after 5522000 ns, '0' after 5522050 ns,
'1' after 5533000 ns, '0' after 5533050 ns,
'1' after 5544000 ns, '0' after 5544050 ns,
'1' after 5555000 ns, '0' after 5555050 ns,
'1' after 5566000 ns, '0' after 5566050 ns,
'1' after 5577000 ns, '0' after 5577050 ns,
'1' after 5588000 ns, '0' after 5588050 ns,
'1' after 5599000 ns, '0' after 5599050 ns,
'1' after 5610000 ns, '0' after 5610050 ns,
'1' after 5621000 ns, '0' after 5621050 ns,
'1' after 5632000 ns, '0' after 5632050 ns,
'1' after 5643000 ns, '0' after 5643050 ns,
'1' after 5654000 ns, '0' after 5654050 ns,
'1' after 5665000 ns, '0' after 5665050 ns,
'1' after 5676000 ns, '0' after 5676050 ns,
'1' after 5687000 ns, '0' after 5687050 ns,
'1' after 5698000 ns, '0' after 5698050 ns,
'1' after 5709000 ns, '0' after 5709050 ns,
'1' after 5720000 ns, '0' after 5720050 ns,
'1' after 5731000 ns, '0' after 5731050 ns,
'1' after 5742000 ns, '0' after 5742050 ns,
'1' after 5753000 ns, '0' after 5753050 ns,
'1' after 5764000 ns, '0' after 5764050 ns,
'1' after 5775000 ns, '0' after 5775050 ns,
'1' after 5786000 ns, '0' after 5786050 ns,
'1' after 5797000 ns, '0' after 5797050 ns,
'1' after 5808000 ns, '0' after 5808050 ns,
'1' after 5819000 ns, '0' after 5819050 ns,
'1' after 5830000 ns, '0' after 5830050 ns,
'1' after 5841000 ns, '0' after 5841050 ns,
'1' after 5852000 ns, '0' after 5852050 ns,
'1' after 5863000 ns, '0' after 5863050 ns,
'1' after 5874000 ns, '0' after 5874050 ns,
'1' after 5885000 ns, '0' after 5885050 ns,
'1' after 5896000 ns, '0' after 5896050 ns,
'1' after 5907000 ns, '0' after 5907050 ns,
'1' after 5918000 ns, '0' after 5918050 ns,
'1' after 5929000 ns, '0' after 5929050 ns,
'1' after 5940000 ns, '0' after 5940050 ns,
'1' after 5951000 ns, '0' after 5951050 ns,
'1' after 5962000 ns, '0' after 5962050 ns,
'1' after 5973000 ns, '0' after 5973050 ns,
'1' after 5984000 ns, '0' after 5984050 ns,
'1' after 5995000 ns, '0' after 5995050 ns,
'1' after 6006000 ns, '0' after 6006050 ns,
'1' after 6017000 ns, '0' after 6017050 ns,
'1' after 6028000 ns, '0' after 6028050 ns,
'1' after 6039000 ns, '0' after 6039050 ns,
'1' after 6050000 ns, '0' after 6050050 ns,
'1' after 6061000 ns, '0' after 6061050 ns,
'1' after 6072000 ns, '0' after 6072050 ns,
'1' after 6083000 ns, '0' after 6083050 ns,
'1' after 6094000 ns, '0' after 6094050 ns,
'1' after 6105000 ns, '0' after 6105050 ns,
'1' after 6116000 ns, '0' after 6116050 ns,
'1' after 6127000 ns, '0' after 6127050 ns,
'1' after 6138000 ns, '0' after 6138050 ns,
'1' after 6149000 ns, '0' after 6149050 ns,
'1' after 6160000 ns, '0' after 6160050 ns,
'1' after 6171000 ns, '0' after 6171050 ns,
'1' after 6182000 ns, '0' after 6182050 ns,
'1' after 6193000 ns, '0' after 6193050 ns,
'1' after 6204000 ns, '0' after 6204050 ns,
'1' after 6215000 ns, '0' after 6215050 ns,
'1' after 6226000 ns, '0' after 6226050 ns,
'1' after 6237000 ns, '0' after 6237050 ns,
'1' after 6248000 ns, '0' after 6248050 ns,
'1' after 6259000 ns, '0' after 6259050 ns,
'1' after 6270000 ns, '0' after 6270050 ns,
'1' after 6281000 ns, '0' after 6281050 ns,
'1' after 6292000 ns, '0' after 6292050 ns,
'1' after 6303000 ns, '0' after 6303050 ns,
'1' after 6314000 ns, '0' after 6314050 ns,
'1' after 6325000 ns, '0' after 6325050 ns,
'1' after 6336000 ns, '0' after 6336050 ns,
'1' after 6347000 ns, '0' after 6347050 ns,
'1' after 6358000 ns, '0' after 6358050 ns,
'1' after 6369000 ns, '0' after 6369050 ns,
'1' after 6380000 ns, '0' after 6380050 ns,
'1' after 6391000 ns, '0' after 6391050 ns,
'1' after 6402000 ns, '0' after 6402050 ns,
'1' after 6413000 ns, '0' after 6413050 ns,
'1' after 6424000 ns, '0' after 6424050 ns,
'1' after 6435000 ns, '0' after 6435050 ns,
'1' after 6446000 ns, '0' after 6446050 ns,
'1' after 6457000 ns, '0' after 6457050 ns,
'1' after 6468000 ns, '0' after 6468050 ns,
'1' after 6479000 ns, '0' after 6479050 ns,
'1' after 6490000 ns, '0' after 6490050 ns,
'1' after 6501000 ns, '0' after 6501050 ns,
'1' after 6512000 ns, '0' after 6512050 ns,
'1' after 6523000 ns, '0' after 6523050 ns,
'1' after 6534000 ns, '0' after 6534050 ns,
'1' after 6545000 ns, '0' after 6545050 ns,
'1' after 6556000 ns, '0' after 6556050 ns,
'1' after 6567000 ns, '0' after 6567050 ns,
'1' after 6578000 ns, '0' after 6578050 ns,
'1' after 6589000 ns, '0' after 6589050 ns,
'1' after 6600000 ns, '0' after 6600050 ns,
'1' after 6611000 ns, '0' after 6611050 ns,
'1' after 6622000 ns, '0' after 6622050 ns,
'1' after 6633000 ns, '0' after 6633050 ns,
'1' after 6644000 ns, '0' after 6644050 ns,
'1' after 6655000 ns, '0' after 6655050 ns,
'1' after 6666000 ns, '0' after 6666050 ns,
'1' after 6677000 ns, '0' after 6677050 ns,
'1' after 6688000 ns, '0' after 6688050 ns,
'1' after 6699000 ns, '0' after 6699050 ns,
'1' after 6710000 ns, '0' after 6710050 ns,
'1' after 6721000 ns, '0' after 6721050 ns,
'1' after 6732000 ns, '0' after 6732050 ns,
'1' after 6743000 ns, '0' after 6743050 ns,
'1' after 6754000 ns, '0' after 6754050 ns,
'1' after 6765000 ns, '0' after 6765050 ns,
'1' after 6776000 ns, '0' after 6776050 ns,
'1' after 6787000 ns, '0' after 6787050 ns,
'1' after 6798000 ns, '0' after 6798050 ns,
'1' after 6809000 ns, '0' after 6809050 ns,
'1' after 6820000 ns, '0' after 6820050 ns,
'1' after 6831000 ns, '0' after 6831050 ns,
'1' after 6842000 ns, '0' after 6842050 ns,
'1' after 6853000 ns, '0' after 6853050 ns,
'1' after 6864000 ns, '0' after 6864050 ns,
'1' after 6875000 ns, '0' after 6875050 ns,
'1' after 6886000 ns, '0' after 6886050 ns,
'1' after 6897000 ns, '0' after 6897050 ns,
'1' after 6908000 ns, '0' after 6908050 ns,
'1' after 6919000 ns, '0' after 6919050 ns,
'1' after 6930000 ns, '0' after 6930050 ns,
'1' after 6941000 ns, '0' after 6941050 ns,
'1' after 6952000 ns, '0' after 6952050 ns,
'1' after 6963000 ns, '0' after 6963050 ns,
'1' after 6974000 ns, '0' after 6974050 ns,
'1' after 6985000 ns, '0' after 6985050 ns,
'1' after 6996000 ns, '0' after 6996050 ns,
'1' after 7007000 ns, '0' after 7007050 ns,
'1' after 7018000 ns, '0' after 7018050 ns,
'1' after 7029000 ns, '0' after 7029050 ns,
'1' after 7040000 ns, '0' after 7040050 ns,
'1' after 7051000 ns, '0' after 7051050 ns,
'1' after 7062000 ns, '0' after 7062050 ns,
'1' after 7073000 ns, '0' after 7073050 ns,
'1' after 7084000 ns, '0' after 7084050 ns,
'1' after 7095000 ns, '0' after 7095050 ns,
'1' after 7106000 ns, '0' after 7106050 ns,
'1' after 7117000 ns, '0' after 7117050 ns,
'1' after 7128000 ns, '0' after 7128050 ns,
'1' after 7139000 ns, '0' after 7139050 ns,
'1' after 7150000 ns, '0' after 7150050 ns,
'1' after 7161000 ns, '0' after 7161050 ns,
'1' after 7172000 ns, '0' after 7172050 ns,
'1' after 7183000 ns, '0' after 7183050 ns,
'1' after 7194000 ns, '0' after 7194050 ns,
'1' after 7205000 ns, '0' after 7205050 ns,
'1' after 7216000 ns, '0' after 7216050 ns,
'1' after 7227000 ns, '0' after 7227050 ns,
'1' after 7238000 ns, '0' after 7238050 ns,
'1' after 7249000 ns, '0' after 7249050 ns,
'1' after 7260000 ns, '0' after 7260050 ns,
'1' after 7271000 ns, '0' after 7271050 ns,
'1' after 7282000 ns, '0' after 7282050 ns,
'1' after 7293000 ns, '0' after 7293050 ns,
'1' after 7304000 ns, '0' after 7304050 ns,
'1' after 7315000 ns, '0' after 7315050 ns,
'1' after 7326000 ns, '0' after 7326050 ns,
'1' after 7337000 ns, '0' after 7337050 ns,
'1' after 7348000 ns, '0' after 7348050 ns,
'1' after 7359000 ns, '0' after 7359050 ns,
'1' after 7370000 ns, '0' after 7370050 ns,
'1' after 7381000 ns, '0' after 7381050 ns,
'1' after 7392000 ns, '0' after 7392050 ns,
'1' after 7403000 ns, '0' after 7403050 ns,
'1' after 7414000 ns, '0' after 7414050 ns,
'1' after 7425000 ns, '0' after 7425050 ns,
'1' after 7436000 ns, '0' after 7436050 ns,
'1' after 7447000 ns, '0' after 7447050 ns,
'1' after 7458000 ns, '0' after 7458050 ns,
'1' after 7469000 ns, '0' after 7469050 ns,
'1' after 7480000 ns, '0' after 7480050 ns,
'1' after 7491000 ns, '0' after 7491050 ns,
'1' after 7502000 ns, '0' after 7502050 ns,
'1' after 7513000 ns, '0' after 7513050 ns,
'1' after 7524000 ns, '0' after 7524050 ns,
'1' after 7535000 ns, '0' after 7535050 ns,
'1' after 7546000 ns, '0' after 7546050 ns,
'1' after 7557000 ns, '0' after 7557050 ns,
'1' after 7568000 ns, '0' after 7568050 ns,
'1' after 7579000 ns, '0' after 7579050 ns,
'1' after 7590000 ns, '0' after 7590050 ns,
'1' after 7601000 ns, '0' after 7601050 ns,
'1' after 7612000 ns, '0' after 7612050 ns,
'1' after 7623000 ns, '0' after 7623050 ns,
'1' after 7634000 ns, '0' after 7634050 ns,
'1' after 7645000 ns, '0' after 7645050 ns,
'1' after 7656000 ns, '0' after 7656050 ns,
'1' after 7667000 ns, '0' after 7667050 ns,
'1' after 7678000 ns, '0' after 7678050 ns,
'1' after 7689000 ns, '0' after 7689050 ns,
'1' after 7700000 ns, '0' after 7700050 ns,
'1' after 7711000 ns, '0' after 7711050 ns,
'1' after 7722000 ns, '0' after 7722050 ns,
'1' after 7733000 ns, '0' after 7733050 ns,
'1' after 7744000 ns, '0' after 7744050 ns,
'1' after 7755000 ns, '0' after 7755050 ns,
'1' after 7766000 ns, '0' after 7766050 ns,
'1' after 7777000 ns, '0' after 7777050 ns,
'1' after 7788000 ns, '0' after 7788050 ns,
'1' after 7799000 ns, '0' after 7799050 ns,
'1' after 7810000 ns, '0' after 7810050 ns,
'1' after 7821000 ns, '0' after 7821050 ns,
'1' after 7832000 ns, '0' after 7832050 ns,
'1' after 7843000 ns, '0' after 7843050 ns,
'1' after 7854000 ns, '0' after 7854050 ns,
'1' after 7865000 ns, '0' after 7865050 ns,
'1' after 7876000 ns, '0' after 7876050 ns,
'1' after 7887000 ns, '0' after 7887050 ns,
'1' after 7898000 ns, '0' after 7898050 ns,
'1' after 7909000 ns, '0' after 7909050 ns,
'1' after 7920000 ns, '0' after 7920050 ns,
'1' after 7931000 ns, '0' after 7931050 ns,
'1' after 7942000 ns, '0' after 7942050 ns,
'1' after 7953000 ns, '0' after 7953050 ns,
'1' after 7964000 ns, '0' after 7964050 ns,
'1' after 7975000 ns, '0' after 7975050 ns,
'1' after 7986000 ns, '0' after 7986050 ns,
'1' after 7997000 ns, '0' after 7997050 ns,
'1' after 8008000 ns, '0' after 8008050 ns,
'1' after 8019000 ns, '0' after 8019050 ns,
'1' after 8030000 ns, '0' after 8030050 ns,
'1' after 8041000 ns, '0' after 8041050 ns,
'1' after 8052000 ns, '0' after 8052050 ns,
'1' after 8063000 ns, '0' after 8063050 ns,
'1' after 8074000 ns, '0' after 8074050 ns,
'1' after 8085000 ns, '0' after 8085050 ns,
'1' after 8096000 ns, '0' after 8096050 ns,
'1' after 8107000 ns, '0' after 8107050 ns,
'1' after 8118000 ns, '0' after 8118050 ns,
'1' after 8129000 ns, '0' after 8129050 ns,
'1' after 8140000 ns, '0' after 8140050 ns,
'1' after 8151000 ns, '0' after 8151050 ns,
'1' after 8162000 ns, '0' after 8162050 ns,
'1' after 8173000 ns, '0' after 8173050 ns,
'1' after 8184000 ns, '0' after 8184050 ns,
'1' after 8195000 ns, '0' after 8195050 ns,
'1' after 8206000 ns, '0' after 8206050 ns,
'1' after 8217000 ns, '0' after 8217050 ns,
'1' after 8228000 ns, '0' after 8228050 ns,
'1' after 8239000 ns, '0' after 8239050 ns,
'1' after 8250000 ns, '0' after 8250050 ns,
'1' after 8261000 ns, '0' after 8261050 ns,
'1' after 8272000 ns, '0' after 8272050 ns,
'1' after 8283000 ns, '0' after 8283050 ns,
'1' after 8294000 ns, '0' after 8294050 ns,
'1' after 8305000 ns, '0' after 8305050 ns,
'1' after 8316000 ns, '0' after 8316050 ns,
'1' after 8327000 ns, '0' after 8327050 ns,
'1' after 8338000 ns, '0' after 8338050 ns,
'1' after 8349000 ns, '0' after 8349050 ns,
'1' after 8360000 ns, '0' after 8360050 ns,
'1' after 8371000 ns, '0' after 8371050 ns,
'1' after 8382000 ns, '0' after 8382050 ns,
'1' after 8393000 ns, '0' after 8393050 ns,
'1' after 8404000 ns, '0' after 8404050 ns,
'1' after 8415000 ns, '0' after 8415050 ns,
'1' after 8426000 ns, '0' after 8426050 ns,
'1' after 8437000 ns, '0' after 8437050 ns,
'1' after 8448000 ns, '0' after 8448050 ns,
'1' after 8459000 ns, '0' after 8459050 ns,
'1' after 8470000 ns, '0' after 8470050 ns,
'1' after 8481000 ns, '0' after 8481050 ns,
'1' after 8492000 ns, '0' after 8492050 ns,
'1' after 8503000 ns, '0' after 8503050 ns,
'1' after 8514000 ns, '0' after 8514050 ns,
'1' after 8525000 ns, '0' after 8525050 ns,
'1' after 8536000 ns, '0' after 8536050 ns,
'1' after 8547000 ns, '0' after 8547050 ns,
'1' after 8558000 ns, '0' after 8558050 ns,
'1' after 8569000 ns, '0' after 8569050 ns,
'1' after 8580000 ns, '0' after 8580050 ns,
'1' after 8591000 ns, '0' after 8591050 ns,
'1' after 8602000 ns, '0' after 8602050 ns,
'1' after 8613000 ns, '0' after 8613050 ns,
'1' after 8624000 ns, '0' after 8624050 ns,
'1' after 8635000 ns, '0' after 8635050 ns,
'1' after 8646000 ns, '0' after 8646050 ns,
'1' after 8657000 ns, '0' after 8657050 ns,
'1' after 8668000 ns, '0' after 8668050 ns,
'1' after 8679000 ns, '0' after 8679050 ns,
'1' after 8690000 ns, '0' after 8690050 ns,
'1' after 8701000 ns, '0' after 8701050 ns,
'1' after 8712000 ns, '0' after 8712050 ns,
'1' after 8723000 ns, '0' after 8723050 ns,
'1' after 8734000 ns, '0' after 8734050 ns,
'1' after 8745000 ns, '0' after 8745050 ns,
'1' after 8756000 ns, '0' after 8756050 ns,
'1' after 8767000 ns, '0' after 8767050 ns,
'1' after 8778000 ns, '0' after 8778050 ns,
'1' after 8789000 ns, '0' after 8789050 ns,
'1' after 8800000 ns, '0' after 8800050 ns,
'1' after 8811000 ns, '0' after 8811050 ns,
'1' after 8822000 ns, '0' after 8822050 ns,
'1' after 8833000 ns, '0' after 8833050 ns,
'1' after 8844000 ns, '0' after 8844050 ns,
'1' after 8855000 ns, '0' after 8855050 ns,
'1' after 8866000 ns, '0' after 8866050 ns,
'1' after 8877000 ns, '0' after 8877050 ns,
'1' after 8888000 ns, '0' after 8888050 ns,
'1' after 8899000 ns, '0' after 8899050 ns,
'1' after 8910000 ns, '0' after 8910050 ns,
'1' after 8921000 ns, '0' after 8921050 ns,
'1' after 8932000 ns, '0' after 8932050 ns,
'1' after 8943000 ns, '0' after 8943050 ns,
'1' after 8954000 ns, '0' after 8954050 ns,
'1' after 8965000 ns, '0' after 8965050 ns,
'1' after 8976000 ns, '0' after 8976050 ns,
'1' after 8987000 ns, '0' after 8987050 ns,
'1' after 8998000 ns, '0' after 8998050 ns,
'1' after 9009000 ns, '0' after 9009050 ns,
'1' after 9020000 ns, '0' after 9020050 ns,
'1' after 9031000 ns, '0' after 9031050 ns,
'1' after 9042000 ns, '0' after 9042050 ns,
'1' after 9053000 ns, '0' after 9053050 ns,
'1' after 9064000 ns, '0' after 9064050 ns,
'1' after 9075000 ns, '0' after 9075050 ns,
'1' after 9086000 ns, '0' after 9086050 ns,
'1' after 9097000 ns, '0' after 9097050 ns,
'1' after 9108000 ns, '0' after 9108050 ns,
'1' after 9119000 ns, '0' after 9119050 ns,
'1' after 9130000 ns, '0' after 9130050 ns,
'1' after 9141000 ns, '0' after 9141050 ns,
'1' after 9152000 ns, '0' after 9152050 ns,
'1' after 9163000 ns, '0' after 9163050 ns,
'1' after 9174000 ns, '0' after 9174050 ns,
'1' after 9185000 ns, '0' after 9185050 ns,
'1' after 9196000 ns, '0' after 9196050 ns,
'1' after 9207000 ns, '0' after 9207050 ns,
'1' after 9218000 ns, '0' after 9218050 ns,
'1' after 9229000 ns, '0' after 9229050 ns,
'1' after 9240000 ns, '0' after 9240050 ns,
'1' after 9251000 ns, '0' after 9251050 ns,
'1' after 9262000 ns, '0' after 9262050 ns,
'1' after 9273000 ns, '0' after 9273050 ns,
'1' after 9284000 ns, '0' after 9284050 ns,
'1' after 9295000 ns, '0' after 9295050 ns,
'1' after 9306000 ns, '0' after 9306050 ns,
'1' after 9317000 ns, '0' after 9317050 ns,
'1' after 9328000 ns, '0' after 9328050 ns,
'1' after 9339000 ns, '0' after 9339050 ns,
'1' after 9350000 ns, '0' after 9350050 ns,
'1' after 9361000 ns, '0' after 9361050 ns,
'1' after 9372000 ns, '0' after 9372050 ns,
'1' after 9383000 ns, '0' after 9383050 ns,
'1' after 9394000 ns, '0' after 9394050 ns,
'1' after 9405000 ns, '0' after 9405050 ns,
'1' after 9416000 ns, '0' after 9416050 ns,
'1' after 9427000 ns, '0' after 9427050 ns,
'1' after 9438000 ns, '0' after 9438050 ns,
'1' after 9449000 ns, '0' after 9449050 ns,
'1' after 9460000 ns, '0' after 9460050 ns,
'1' after 9471000 ns, '0' after 9471050 ns,
'1' after 9482000 ns, '0' after 9482050 ns,
'1' after 9493000 ns, '0' after 9493050 ns,
'1' after 9504000 ns, '0' after 9504050 ns,
'1' after 9515000 ns, '0' after 9515050 ns,
'1' after 9526000 ns, '0' after 9526050 ns,
'1' after 9537000 ns, '0' after 9537050 ns,
'1' after 9548000 ns, '0' after 9548050 ns,
'1' after 9559000 ns, '0' after 9559050 ns,
'1' after 9570000 ns, '0' after 9570050 ns,
'1' after 9581000 ns, '0' after 9581050 ns,
'1' after 9592000 ns, '0' after 9592050 ns,
'1' after 9603000 ns, '0' after 9603050 ns,
'1' after 9614000 ns, '0' after 9614050 ns,
'1' after 9625000 ns, '0' after 9625050 ns,
'1' after 9636000 ns, '0' after 9636050 ns,
'1' after 9647000 ns, '0' after 9647050 ns,
'1' after 9658000 ns, '0' after 9658050 ns,
'1' after 9669000 ns, '0' after 9669050 ns,
'1' after 9680000 ns, '0' after 9680050 ns,
'1' after 9691000 ns, '0' after 9691050 ns,
'1' after 9702000 ns, '0' after 9702050 ns,
'1' after 9713000 ns, '0' after 9713050 ns,
'1' after 9724000 ns, '0' after 9724050 ns,
'1' after 9735000 ns, '0' after 9735050 ns,
'1' after 9746000 ns, '0' after 9746050 ns,
'1' after 9757000 ns, '0' after 9757050 ns,
'1' after 9768000 ns, '0' after 9768050 ns,
'1' after 9779000 ns, '0' after 9779050 ns,
'1' after 9790000 ns, '0' after 9790050 ns,
'1' after 9801000 ns, '0' after 9801050 ns,
'1' after 9812000 ns, '0' after 9812050 ns,
'1' after 9823000 ns, '0' after 9823050 ns,
'1' after 9834000 ns, '0' after 9834050 ns,
'1' after 9845000 ns, '0' after 9845050 ns,
'1' after 9856000 ns, '0' after 9856050 ns,
'1' after 9867000 ns, '0' after 9867050 ns,
'1' after 9878000 ns, '0' after 9878050 ns,
'1' after 9889000 ns, '0' after 9889050 ns,
'1' after 9900000 ns, '0' after 9900050 ns,
'1' after 9911000 ns, '0' after 9911050 ns,
'1' after 9922000 ns, '0' after 9922050 ns,
'1' after 9933000 ns, '0' after 9933050 ns,
'1' after 9944000 ns, '0' after 9944050 ns,
'1' after 9955000 ns, '0' after 9955050 ns,
'1' after 9966000 ns, '0' after 9966050 ns,
'1' after 9977000 ns, '0' after 9977050 ns,
'1' after 9988000 ns, '0' after 9988050 ns,
'1' after 9999000 ns, '0' after 9999050 ns,
'1' after 10010000 ns, '0' after 10010050 ns,
'1' after 10021000 ns, '0' after 10021050 ns,
'1' after 10032000 ns, '0' after 10032050 ns,
'1' after 10043000 ns, '0' after 10043050 ns,
'1' after 10054000 ns, '0' after 10054050 ns,
'1' after 10065000 ns, '0' after 10065050 ns,
'1' after 10076000 ns, '0' after 10076050 ns,
'1' after 10087000 ns, '0' after 10087050 ns,
'1' after 10098000 ns, '0' after 10098050 ns,
'1' after 10109000 ns, '0' after 10109050 ns,
'1' after 10120000 ns, '0' after 10120050 ns,
'1' after 10131000 ns, '0' after 10131050 ns,
'1' after 10142000 ns, '0' after 10142050 ns,
'1' after 10153000 ns, '0' after 10153050 ns,
'1' after 10164000 ns, '0' after 10164050 ns,
'1' after 10175000 ns, '0' after 10175050 ns,
'1' after 10186000 ns, '0' after 10186050 ns,
'1' after 10197000 ns, '0' after 10197050 ns,
'1' after 10208000 ns, '0' after 10208050 ns,
'1' after 10219000 ns, '0' after 10219050 ns,
'1' after 10230000 ns, '0' after 10230050 ns,
'1' after 10241000 ns, '0' after 10241050 ns,
'1' after 10252000 ns, '0' after 10252050 ns,
'1' after 10263000 ns, '0' after 10263050 ns,
'1' after 10274000 ns, '0' after 10274050 ns,
'1' after 10285000 ns, '0' after 10285050 ns,
'1' after 10296000 ns, '0' after 10296050 ns,
'1' after 10307000 ns, '0' after 10307050 ns,
'1' after 10318000 ns, '0' after 10318050 ns,
'1' after 10329000 ns, '0' after 10329050 ns,
'1' after 10340000 ns, '0' after 10340050 ns,
'1' after 10351000 ns, '0' after 10351050 ns,
'1' after 10362000 ns, '0' after 10362050 ns,
'1' after 10373000 ns, '0' after 10373050 ns,
'1' after 10384000 ns, '0' after 10384050 ns,
'1' after 10395000 ns, '0' after 10395050 ns,
'1' after 10406000 ns, '0' after 10406050 ns,
'1' after 10417000 ns, '0' after 10417050 ns,
'1' after 10428000 ns, '0' after 10428050 ns,
'1' after 10439000 ns, '0' after 10439050 ns,
'1' after 10450000 ns, '0' after 10450050 ns,
'1' after 10461000 ns, '0' after 10461050 ns,
'1' after 10472000 ns, '0' after 10472050 ns,
'1' after 10483000 ns, '0' after 10483050 ns,
'1' after 10494000 ns, '0' after 10494050 ns,
'1' after 10505000 ns, '0' after 10505050 ns,
'1' after 10516000 ns, '0' after 10516050 ns,
'1' after 10527000 ns, '0' after 10527050 ns,
'1' after 10538000 ns, '0' after 10538050 ns,
'1' after 10549000 ns, '0' after 10549050 ns,
'1' after 10560000 ns, '0' after 10560050 ns,
'1' after 10571000 ns, '0' after 10571050 ns,
'1' after 10582000 ns, '0' after 10582050 ns,
'1' after 10593000 ns, '0' after 10593050 ns,
'1' after 10604000 ns, '0' after 10604050 ns,
'1' after 10615000 ns, '0' after 10615050 ns,
'1' after 10626000 ns, '0' after 10626050 ns,
'1' after 10637000 ns, '0' after 10637050 ns,
'1' after 10648000 ns, '0' after 10648050 ns,
'1' after 10659000 ns, '0' after 10659050 ns,
'1' after 10670000 ns, '0' after 10670050 ns,
'1' after 10681000 ns, '0' after 10681050 ns,
'1' after 10692000 ns, '0' after 10692050 ns,
'1' after 10703000 ns, '0' after 10703050 ns,
'1' after 10714000 ns, '0' after 10714050 ns,
'1' after 10725000 ns, '0' after 10725050 ns,
'1' after 10736000 ns, '0' after 10736050 ns,
'1' after 10747000 ns, '0' after 10747050 ns,
'1' after 10758000 ns, '0' after 10758050 ns,
'1' after 10769000 ns, '0' after 10769050 ns,
'1' after 10780000 ns, '0' after 10780050 ns,
'1' after 10791000 ns, '0' after 10791050 ns,
'1' after 10802000 ns, '0' after 10802050 ns,
'1' after 10813000 ns, '0' after 10813050 ns,
'1' after 10824000 ns, '0' after 10824050 ns,
'1' after 10835000 ns, '0' after 10835050 ns,
'1' after 10846000 ns, '0' after 10846050 ns,
'1' after 10857000 ns, '0' after 10857050 ns,
'1' after 10868000 ns, '0' after 10868050 ns,
'1' after 10879000 ns, '0' after 10879050 ns,
'1' after 10890000 ns, '0' after 10890050 ns,
'1' after 10901000 ns, '0' after 10901050 ns,
'1' after 10912000 ns, '0' after 10912050 ns,
'1' after 10923000 ns, '0' after 10923050 ns,
'1' after 10934000 ns, '0' after 10934050 ns,
'1' after 10945000 ns, '0' after 10945050 ns,
'1' after 10956000 ns, '0' after 10956050 ns,
'1' after 10967000 ns, '0' after 10967050 ns,
'1' after 10978000 ns, '0' after 10978050 ns,
'1' after 10989000 ns, '0' after 10989050 ns,
'1' after 11000000 ns, '0' after 11000050 ns,
'1' after 11011000 ns, '0' after 11011050 ns,
'1' after 11022000 ns, '0' after 11022050 ns,
'1' after 11033000 ns, '0' after 11033050 ns,
'1' after 11044000 ns, '0' after 11044050 ns,
'1' after 11055000 ns, '0' after 11055050 ns,
'1' after 11066000 ns, '0' after 11066050 ns,
'1' after 11077000 ns, '0' after 11077050 ns,
'1' after 11088000 ns, '0' after 11088050 ns,
'1' after 11099000 ns, '0' after 11099050 ns,
'1' after 11110000 ns, '0' after 11110050 ns,
'1' after 11121000 ns, '0' after 11121050 ns,
'1' after 11132000 ns, '0' after 11132050 ns,
'1' after 11143000 ns, '0' after 11143050 ns,
'1' after 11154000 ns, '0' after 11154050 ns,
'1' after 11165000 ns, '0' after 11165050 ns,
'1' after 11176000 ns, '0' after 11176050 ns,
'1' after 11187000 ns, '0' after 11187050 ns,
'1' after 11198000 ns, '0' after 11198050 ns,
'1' after 11209000 ns, '0' after 11209050 ns,
'1' after 11220000 ns, '0' after 11220050 ns,
'1' after 11231000 ns, '0' after 11231050 ns,
'1' after 11242000 ns, '0' after 11242050 ns,
'1' after 11253000 ns, '0' after 11253050 ns,
'1' after 11264000 ns, '0' after 11264050 ns,
'1' after 11275000 ns, '0' after 11275050 ns,
'1' after 11286000 ns, '0' after 11286050 ns,
'1' after 11297000 ns, '0' after 11297050 ns,
'1' after 11308000 ns, '0' after 11308050 ns,
'1' after 11319000 ns, '0' after 11319050 ns,
'1' after 11330000 ns, '0' after 11330050 ns,
'1' after 11341000 ns, '0' after 11341050 ns,
'1' after 11352000 ns, '0' after 11352050 ns,
'1' after 11363000 ns, '0' after 11363050 ns,
'1' after 11374000 ns, '0' after 11374050 ns,
'1' after 11385000 ns, '0' after 11385050 ns,
'1' after 11396000 ns, '0' after 11396050 ns,
'1' after 11407000 ns, '0' after 11407050 ns,
'1' after 11418000 ns, '0' after 11418050 ns,
'1' after 11429000 ns, '0' after 11429050 ns,
'1' after 11440000 ns, '0' after 11440050 ns,
'1' after 11451000 ns, '0' after 11451050 ns,
'1' after 11462000 ns, '0' after 11462050 ns,
'1' after 11473000 ns, '0' after 11473050 ns,
'1' after 11484000 ns, '0' after 11484050 ns,
'1' after 11495000 ns, '0' after 11495050 ns,
'1' after 11506000 ns, '0' after 11506050 ns,
'1' after 11517000 ns, '0' after 11517050 ns,
'1' after 11528000 ns, '0' after 11528050 ns,
'1' after 11539000 ns, '0' after 11539050 ns,
'1' after 11550000 ns, '0' after 11550050 ns,
'1' after 11561000 ns, '0' after 11561050 ns,
'1' after 11572000 ns, '0' after 11572050 ns,
'1' after 11583000 ns, '0' after 11583050 ns,
'1' after 11594000 ns, '0' after 11594050 ns,
'1' after 11605000 ns, '0' after 11605050 ns,
'1' after 11616000 ns, '0' after 11616050 ns,
'1' after 11627000 ns, '0' after 11627050 ns,
'1' after 11638000 ns, '0' after 11638050 ns,
'1' after 11649000 ns, '0' after 11649050 ns,
'1' after 11660000 ns, '0' after 11660050 ns,
'1' after 11671000 ns, '0' after 11671050 ns,
'1' after 11682000 ns, '0' after 11682050 ns,
'1' after 11693000 ns, '0' after 11693050 ns,
'1' after 11704000 ns, '0' after 11704050 ns,
'1' after 11715000 ns, '0' after 11715050 ns,
'1' after 11726000 ns, '0' after 11726050 ns,
'1' after 11737000 ns, '0' after 11737050 ns,
'1' after 11748000 ns, '0' after 11748050 ns,
'1' after 11759000 ns, '0' after 11759050 ns,
'1' after 11770000 ns, '0' after 11770050 ns,
'1' after 11781000 ns, '0' after 11781050 ns,
'1' after 11792000 ns, '0' after 11792050 ns,
'1' after 11803000 ns, '0' after 11803050 ns,
'1' after 11814000 ns, '0' after 11814050 ns,
'1' after 11825000 ns, '0' after 11825050 ns,
'1' after 11836000 ns, '0' after 11836050 ns,
'1' after 11847000 ns, '0' after 11847050 ns,
'1' after 11858000 ns, '0' after 11858050 ns,
'1' after 11869000 ns, '0' after 11869050 ns,
'1' after 11880000 ns, '0' after 11880050 ns,
'1' after 11891000 ns, '0' after 11891050 ns,
'1' after 11902000 ns, '0' after 11902050 ns,
'1' after 11913000 ns, '0' after 11913050 ns,
'1' after 11924000 ns, '0' after 11924050 ns,
'1' after 11935000 ns, '0' after 11935050 ns,
'1' after 11946000 ns, '0' after 11946050 ns,
'1' after 11957000 ns, '0' after 11957050 ns,
'1' after 11968000 ns, '0' after 11968050 ns,
'1' after 11979000 ns, '0' after 11979050 ns,
'1' after 11990000 ns, '0' after 11990050 ns,
'1' after 12001000 ns, '0' after 12001050 ns,
'1' after 12012000 ns, '0' after 12012050 ns,
'1' after 12023000 ns, '0' after 12023050 ns,
'1' after 12034000 ns, '0' after 12034050 ns,
'1' after 12045000 ns, '0' after 12045050 ns,
'1' after 12056000 ns, '0' after 12056050 ns,
'1' after 12067000 ns, '0' after 12067050 ns,
'1' after 12078000 ns, '0' after 12078050 ns,
'1' after 12089000 ns, '0' after 12089050 ns,
'1' after 12100000 ns, '0' after 12100050 ns,
'1' after 12111000 ns, '0' after 12111050 ns,
'1' after 12122000 ns, '0' after 12122050 ns,
'1' after 12133000 ns, '0' after 12133050 ns,
'1' after 12144000 ns, '0' after 12144050 ns,
'1' after 12155000 ns, '0' after 12155050 ns,
'1' after 12166000 ns, '0' after 12166050 ns,
'1' after 12177000 ns, '0' after 12177050 ns,
'1' after 12188000 ns, '0' after 12188050 ns,
'1' after 12199000 ns, '0' after 12199050 ns,
'1' after 12210000 ns, '0' after 12210050 ns,
'1' after 12221000 ns, '0' after 12221050 ns,
'1' after 12232000 ns, '0' after 12232050 ns,
'1' after 12243000 ns, '0' after 12243050 ns,
'1' after 12254000 ns, '0' after 12254050 ns,
'1' after 12265000 ns, '0' after 12265050 ns,
'1' after 12276000 ns, '0' after 12276050 ns,
'1' after 12287000 ns, '0' after 12287050 ns,
'1' after 12298000 ns, '0' after 12298050 ns,
'1' after 12309000 ns, '0' after 12309050 ns,
'1' after 12320000 ns, '0' after 12320050 ns,
'1' after 12331000 ns, '0' after 12331050 ns,
'1' after 12342000 ns, '0' after 12342050 ns,
'1' after 12353000 ns, '0' after 12353050 ns,
'1' after 12364000 ns, '0' after 12364050 ns,
'1' after 12375000 ns, '0' after 12375050 ns,
'1' after 12386000 ns, '0' after 12386050 ns,
'1' after 12397000 ns, '0' after 12397050 ns,
'1' after 12408000 ns, '0' after 12408050 ns,
'1' after 12419000 ns, '0' after 12419050 ns,
'1' after 12430000 ns, '0' after 12430050 ns,
'1' after 12441000 ns, '0' after 12441050 ns,
'1' after 12452000 ns, '0' after 12452050 ns,
'1' after 12463000 ns, '0' after 12463050 ns,
'1' after 12474000 ns, '0' after 12474050 ns,
'1' after 12485000 ns, '0' after 12485050 ns,
'1' after 12496000 ns, '0' after 12496050 ns,
'1' after 12507000 ns, '0' after 12507050 ns,
'1' after 12518000 ns, '0' after 12518050 ns,
'1' after 12529000 ns, '0' after 12529050 ns,
'1' after 12540000 ns, '0' after 12540050 ns,
'1' after 12551000 ns, '0' after 12551050 ns,
'1' after 12562000 ns, '0' after 12562050 ns,
'1' after 12573000 ns, '0' after 12573050 ns,
'1' after 12584000 ns, '0' after 12584050 ns,
'1' after 12595000 ns, '0' after 12595050 ns,
'1' after 12606000 ns, '0' after 12606050 ns,
'1' after 12617000 ns, '0' after 12617050 ns,
'1' after 12628000 ns, '0' after 12628050 ns,
'1' after 12639000 ns, '0' after 12639050 ns,
'1' after 12650000 ns, '0' after 12650050 ns,
'1' after 12661000 ns, '0' after 12661050 ns,
'1' after 12672000 ns, '0' after 12672050 ns,
'1' after 12683000 ns, '0' after 12683050 ns,
'1' after 12694000 ns, '0' after 12694050 ns,
'1' after 12705000 ns, '0' after 12705050 ns,
'1' after 12716000 ns, '0' after 12716050 ns,
'1' after 12727000 ns, '0' after 12727050 ns,
'1' after 12738000 ns, '0' after 12738050 ns,
'1' after 12749000 ns, '0' after 12749050 ns,
'1' after 12760000 ns, '0' after 12760050 ns,
'1' after 12771000 ns, '0' after 12771050 ns,
'1' after 12782000 ns, '0' after 12782050 ns,
'1' after 12793000 ns, '0' after 12793050 ns,
'1' after 12804000 ns, '0' after 12804050 ns,
'1' after 12815000 ns, '0' after 12815050 ns,
'1' after 12826000 ns, '0' after 12826050 ns,
'1' after 12837000 ns, '0' after 12837050 ns,
'1' after 12848000 ns, '0' after 12848050 ns,
'1' after 12859000 ns, '0' after 12859050 ns,
'1' after 12870000 ns, '0' after 12870050 ns,
'1' after 12881000 ns, '0' after 12881050 ns,
'1' after 12892000 ns, '0' after 12892050 ns,
'1' after 12903000 ns, '0' after 12903050 ns,
'1' after 12914000 ns, '0' after 12914050 ns,
'1' after 12925000 ns, '0' after 12925050 ns,
'1' after 12936000 ns, '0' after 12936050 ns,
'1' after 12947000 ns, '0' after 12947050 ns,
'1' after 12958000 ns, '0' after 12958050 ns,
'1' after 12969000 ns, '0' after 12969050 ns,
'1' after 12980000 ns, '0' after 12980050 ns,
'1' after 12991000 ns, '0' after 12991050 ns,
'1' after 13002000 ns, '0' after 13002050 ns,
'1' after 13013000 ns, '0' after 13013050 ns,
'1' after 13024000 ns, '0' after 13024050 ns,
'1' after 13035000 ns, '0' after 13035050 ns,
'1' after 13046000 ns, '0' after 13046050 ns,
'1' after 13057000 ns, '0' after 13057050 ns,
'1' after 13068000 ns, '0' after 13068050 ns,
'1' after 13079000 ns, '0' after 13079050 ns,
'1' after 13090000 ns, '0' after 13090050 ns,
'1' after 13101000 ns, '0' after 13101050 ns,
'1' after 13112000 ns, '0' after 13112050 ns,
'1' after 13123000 ns, '0' after 13123050 ns,
'1' after 13134000 ns, '0' after 13134050 ns,
'1' after 13145000 ns, '0' after 13145050 ns,
'1' after 13156000 ns, '0' after 13156050 ns,
'1' after 13167000 ns, '0' after 13167050 ns,
'1' after 13178000 ns, '0' after 13178050 ns,
'1' after 13189000 ns, '0' after 13189050 ns,
'1' after 13200000 ns, '0' after 13200050 ns,
'1' after 13211000 ns, '0' after 13211050 ns,
'1' after 13222000 ns, '0' after 13222050 ns,
'1' after 13233000 ns, '0' after 13233050 ns,
'1' after 13244000 ns, '0' after 13244050 ns,
'1' after 13255000 ns, '0' after 13255050 ns,
'1' after 13266000 ns, '0' after 13266050 ns,
'1' after 13277000 ns, '0' after 13277050 ns,
'1' after 13288000 ns, '0' after 13288050 ns,
'1' after 13299000 ns, '0' after 13299050 ns,
'1' after 13310000 ns, '0' after 13310050 ns,
'1' after 13321000 ns, '0' after 13321050 ns,
'1' after 13332000 ns, '0' after 13332050 ns,
'1' after 13343000 ns, '0' after 13343050 ns,
'1' after 13354000 ns, '0' after 13354050 ns,
'1' after 13365000 ns, '0' after 13365050 ns,
'1' after 13376000 ns, '0' after 13376050 ns,
'1' after 13387000 ns, '0' after 13387050 ns,
'1' after 13398000 ns, '0' after 13398050 ns,
'1' after 13409000 ns, '0' after 13409050 ns,
'1' after 13420000 ns, '0' after 13420050 ns,
'1' after 13431000 ns, '0' after 13431050 ns,
'1' after 13442000 ns, '0' after 13442050 ns,
'1' after 13453000 ns, '0' after 13453050 ns,
'1' after 13464000 ns, '0' after 13464050 ns,
'1' after 13475000 ns, '0' after 13475050 ns,
'1' after 13486000 ns, '0' after 13486050 ns,
'1' after 13497000 ns, '0' after 13497050 ns,
'1' after 13508000 ns, '0' after 13508050 ns,
'1' after 13519000 ns, '0' after 13519050 ns,
'1' after 13530000 ns, '0' after 13530050 ns,
'1' after 13541000 ns, '0' after 13541050 ns,
'1' after 13552000 ns, '0' after 13552050 ns,
'1' after 13563000 ns, '0' after 13563050 ns,
'1' after 13574000 ns, '0' after 13574050 ns,
'1' after 13585000 ns, '0' after 13585050 ns,
'1' after 13596000 ns, '0' after 13596050 ns,
'1' after 13607000 ns, '0' after 13607050 ns,
'1' after 13618000 ns, '0' after 13618050 ns,
'1' after 13629000 ns, '0' after 13629050 ns,
'1' after 13640000 ns, '0' after 13640050 ns,
'1' after 13651000 ns, '0' after 13651050 ns,
'1' after 13662000 ns, '0' after 13662050 ns,
'1' after 13673000 ns, '0' after 13673050 ns,
'1' after 13684000 ns, '0' after 13684050 ns,
'1' after 13695000 ns, '0' after 13695050 ns,
'1' after 13706000 ns, '0' after 13706050 ns,
'1' after 13717000 ns, '0' after 13717050 ns,
'1' after 13728000 ns, '0' after 13728050 ns,
'1' after 13739000 ns, '0' after 13739050 ns,
'1' after 13750000 ns, '0' after 13750050 ns,
'1' after 13761000 ns, '0' after 13761050 ns,
'1' after 13772000 ns, '0' after 13772050 ns,
'1' after 13783000 ns, '0' after 13783050 ns,
'1' after 13794000 ns, '0' after 13794050 ns,
'1' after 13805000 ns, '0' after 13805050 ns,
'1' after 13816000 ns, '0' after 13816050 ns,
'1' after 13827000 ns, '0' after 13827050 ns,
'1' after 13838000 ns, '0' after 13838050 ns,
'1' after 13849000 ns, '0' after 13849050 ns,
'1' after 13860000 ns, '0' after 13860050 ns,
'1' after 13871000 ns, '0' after 13871050 ns,
'1' after 13882000 ns, '0' after 13882050 ns,
'1' after 13893000 ns, '0' after 13893050 ns,
'1' after 13904000 ns, '0' after 13904050 ns,
'1' after 13915000 ns, '0' after 13915050 ns,
'1' after 13926000 ns, '0' after 13926050 ns,
'1' after 13937000 ns, '0' after 13937050 ns,
'1' after 13948000 ns, '0' after 13948050 ns,
'1' after 13959000 ns, '0' after 13959050 ns,
'1' after 13970000 ns, '0' after 13970050 ns,
'1' after 13981000 ns, '0' after 13981050 ns,
'1' after 13992000 ns, '0' after 13992050 ns,
'1' after 14003000 ns, '0' after 14003050 ns,
'1' after 14014000 ns, '0' after 14014050 ns,
'1' after 14025000 ns, '0' after 14025050 ns,
'1' after 14036000 ns, '0' after 14036050 ns,
'1' after 14047000 ns, '0' after 14047050 ns,
'1' after 14058000 ns, '0' after 14058050 ns,
'1' after 14069000 ns, '0' after 14069050 ns,
'1' after 14080000 ns, '0' after 14080050 ns,
'1' after 14091000 ns, '0' after 14091050 ns,
'1' after 14102000 ns, '0' after 14102050 ns,
'1' after 14113000 ns, '0' after 14113050 ns,
'1' after 14124000 ns, '0' after 14124050 ns,
'1' after 14135000 ns, '0' after 14135050 ns,
'1' after 14146000 ns, '0' after 14146050 ns,
'1' after 14157000 ns, '0' after 14157050 ns,
'1' after 14168000 ns, '0' after 14168050 ns,
'1' after 14179000 ns, '0' after 14179050 ns,
'1' after 14190000 ns, '0' after 14190050 ns,
'1' after 14201000 ns, '0' after 14201050 ns,
'1' after 14212000 ns, '0' after 14212050 ns,
'1' after 14223000 ns, '0' after 14223050 ns,
'1' after 14234000 ns, '0' after 14234050 ns,
'1' after 14245000 ns, '0' after 14245050 ns,
'1' after 14256000 ns, '0' after 14256050 ns,
'1' after 14267000 ns, '0' after 14267050 ns,
'1' after 14278000 ns, '0' after 14278050 ns,
'1' after 14289000 ns, '0' after 14289050 ns,
'1' after 14300000 ns, '0' after 14300050 ns,
'1' after 14311000 ns, '0' after 14311050 ns,
'1' after 14322000 ns, '0' after 14322050 ns,
'1' after 14333000 ns, '0' after 14333050 ns,
'1' after 14344000 ns, '0' after 14344050 ns,
'1' after 14355000 ns, '0' after 14355050 ns,
'1' after 14366000 ns, '0' after 14366050 ns,
'1' after 14377000 ns, '0' after 14377050 ns,
'1' after 14388000 ns, '0' after 14388050 ns,
'1' after 14399000 ns, '0' after 14399050 ns,
'1' after 14410000 ns, '0' after 14410050 ns,
'1' after 14421000 ns, '0' after 14421050 ns,
'1' after 14432000 ns, '0' after 14432050 ns,
'1' after 14443000 ns, '0' after 14443050 ns,
'1' after 14454000 ns, '0' after 14454050 ns,
'1' after 14465000 ns, '0' after 14465050 ns,
'1' after 14476000 ns, '0' after 14476050 ns,
'1' after 14487000 ns, '0' after 14487050 ns,
'1' after 14498000 ns, '0' after 14498050 ns,
'1' after 14509000 ns, '0' after 14509050 ns,
'1' after 14520000 ns, '0' after 14520050 ns,
'1' after 14531000 ns, '0' after 14531050 ns,
'1' after 14542000 ns, '0' after 14542050 ns,
'1' after 14553000 ns, '0' after 14553050 ns,
'1' after 14564000 ns, '0' after 14564050 ns,
'1' after 14575000 ns, '0' after 14575050 ns,
'1' after 14586000 ns, '0' after 14586050 ns,
'1' after 14597000 ns, '0' after 14597050 ns,
'1' after 14608000 ns, '0' after 14608050 ns,
'1' after 14619000 ns, '0' after 14619050 ns,
'1' after 14630000 ns, '0' after 14630050 ns,
'1' after 14641000 ns, '0' after 14641050 ns,
'1' after 14652000 ns, '0' after 14652050 ns,
'1' after 14663000 ns, '0' after 14663050 ns,
'1' after 14674000 ns, '0' after 14674050 ns,
'1' after 14685000 ns, '0' after 14685050 ns,
'1' after 14696000 ns, '0' after 14696050 ns,
'1' after 14707000 ns, '0' after 14707050 ns,
'1' after 14718000 ns, '0' after 14718050 ns,
'1' after 14729000 ns, '0' after 14729050 ns,
'1' after 14740000 ns, '0' after 14740050 ns,
'1' after 14751000 ns, '0' after 14751050 ns,
'1' after 14762000 ns, '0' after 14762050 ns,
'1' after 14773000 ns, '0' after 14773050 ns,
'1' after 14784000 ns, '0' after 14784050 ns,
'1' after 14795000 ns, '0' after 14795050 ns,
'1' after 14806000 ns, '0' after 14806050 ns,
'1' after 14817000 ns, '0' after 14817050 ns,
'1' after 14828000 ns, '0' after 14828050 ns,
'1' after 14839000 ns, '0' after 14839050 ns,
'1' after 14850000 ns, '0' after 14850050 ns,
'1' after 14861000 ns, '0' after 14861050 ns,
'1' after 14872000 ns, '0' after 14872050 ns,
'1' after 14883000 ns, '0' after 14883050 ns,
'1' after 14894000 ns, '0' after 14894050 ns,
'1' after 14905000 ns, '0' after 14905050 ns,
'1' after 14916000 ns, '0' after 14916050 ns,
'1' after 14927000 ns, '0' after 14927050 ns,
'1' after 14938000 ns, '0' after 14938050 ns,
'1' after 14949000 ns, '0' after 14949050 ns,
'1' after 14960000 ns, '0' after 14960050 ns,
'1' after 14971000 ns, '0' after 14971050 ns,
'1' after 14982000 ns, '0' after 14982050 ns,
'1' after 14993000 ns, '0' after 14993050 ns,
'1' after 15004000 ns, '0' after 15004050 ns,
'1' after 15015000 ns, '0' after 15015050 ns,
'1' after 15026000 ns, '0' after 15026050 ns,
'1' after 15037000 ns, '0' after 15037050 ns,
'1' after 15048000 ns, '0' after 15048050 ns,
'1' after 15059000 ns, '0' after 15059050 ns,
'1' after 15070000 ns, '0' after 15070050 ns,
'1' after 15081000 ns, '0' after 15081050 ns,
'1' after 15092000 ns, '0' after 15092050 ns,
'1' after 15103000 ns, '0' after 15103050 ns,
'1' after 15114000 ns, '0' after 15114050 ns,
'1' after 15125000 ns, '0' after 15125050 ns,
'1' after 15136000 ns, '0' after 15136050 ns,
'1' after 15147000 ns, '0' after 15147050 ns,
'1' after 15158000 ns, '0' after 15158050 ns,
'1' after 15169000 ns, '0' after 15169050 ns,
'1' after 15180000 ns, '0' after 15180050 ns,
'1' after 15191000 ns, '0' after 15191050 ns,
'1' after 15202000 ns, '0' after 15202050 ns,
'1' after 15213000 ns, '0' after 15213050 ns,
'1' after 15224000 ns, '0' after 15224050 ns,
'1' after 15235000 ns, '0' after 15235050 ns,
'1' after 15246000 ns, '0' after 15246050 ns,
'1' after 15257000 ns, '0' after 15257050 ns,
'1' after 15268000 ns, '0' after 15268050 ns,
'1' after 15279000 ns, '0' after 15279050 ns,
'1' after 15290000 ns, '0' after 15290050 ns,
'1' after 15301000 ns, '0' after 15301050 ns,
'1' after 15312000 ns, '0' after 15312050 ns,
'1' after 15323000 ns, '0' after 15323050 ns,
'1' after 15334000 ns, '0' after 15334050 ns,
'1' after 15345000 ns, '0' after 15345050 ns,
'1' after 15356000 ns, '0' after 15356050 ns,
'1' after 15367000 ns, '0' after 15367050 ns,
'1' after 15378000 ns, '0' after 15378050 ns,
'1' after 15389000 ns, '0' after 15389050 ns,
'1' after 15400000 ns, '0' after 15400050 ns,
'1' after 15411000 ns, '0' after 15411050 ns,
'1' after 15422000 ns, '0' after 15422050 ns,
'1' after 15433000 ns, '0' after 15433050 ns,
'1' after 15444000 ns, '0' after 15444050 ns,
'1' after 15455000 ns, '0' after 15455050 ns,
'1' after 15466000 ns, '0' after 15466050 ns,
'1' after 15477000 ns, '0' after 15477050 ns,
'1' after 15488000 ns, '0' after 15488050 ns,
'1' after 15499000 ns, '0' after 15499050 ns,
'1' after 15510000 ns, '0' after 15510050 ns,
'1' after 15521000 ns, '0' after 15521050 ns,
'1' after 15532000 ns, '0' after 15532050 ns,
'1' after 15543000 ns, '0' after 15543050 ns,
'1' after 15554000 ns, '0' after 15554050 ns,
'1' after 15565000 ns, '0' after 15565050 ns,
'1' after 15576000 ns, '0' after 15576050 ns,
'1' after 15587000 ns, '0' after 15587050 ns,
'1' after 15598000 ns, '0' after 15598050 ns,
'1' after 15609000 ns, '0' after 15609050 ns,
'1' after 15620000 ns, '0' after 15620050 ns,
'1' after 15631000 ns, '0' after 15631050 ns,
'1' after 15642000 ns, '0' after 15642050 ns,
'1' after 15653000 ns, '0' after 15653050 ns,
'1' after 15664000 ns, '0' after 15664050 ns,
'1' after 15675000 ns, '0' after 15675050 ns,
'1' after 15686000 ns, '0' after 15686050 ns,
'1' after 15697000 ns, '0' after 15697050 ns,
'1' after 15708000 ns, '0' after 15708050 ns,
'1' after 15719000 ns, '0' after 15719050 ns,
'1' after 15730000 ns, '0' after 15730050 ns,
'1' after 15741000 ns, '0' after 15741050 ns,
'1' after 15752000 ns, '0' after 15752050 ns,
'1' after 15763000 ns, '0' after 15763050 ns,
'1' after 15774000 ns, '0' after 15774050 ns,
'1' after 15785000 ns, '0' after 15785050 ns,
'1' after 15796000 ns, '0' after 15796050 ns,
'1' after 15807000 ns, '0' after 15807050 ns,
'1' after 15818000 ns, '0' after 15818050 ns,
'1' after 15829000 ns, '0' after 15829050 ns,
'1' after 15840000 ns, '0' after 15840050 ns,
'1' after 15851000 ns, '0' after 15851050 ns,
'1' after 15862000 ns, '0' after 15862050 ns,
'1' after 15873000 ns, '0' after 15873050 ns,
'1' after 15884000 ns, '0' after 15884050 ns,
'1' after 15895000 ns, '0' after 15895050 ns,
'1' after 15906000 ns, '0' after 15906050 ns,
'1' after 15917000 ns, '0' after 15917050 ns,
'1' after 15928000 ns, '0' after 15928050 ns,
'1' after 15939000 ns, '0' after 15939050 ns,
'1' after 15950000 ns, '0' after 15950050 ns,
'1' after 15961000 ns, '0' after 15961050 ns,
'1' after 15972000 ns, '0' after 15972050 ns,
'1' after 15983000 ns, '0' after 15983050 ns,
'1' after 15994000 ns, '0' after 15994050 ns,
'1' after 16005000 ns, '0' after 16005050 ns,
'1' after 16016000 ns, '0' after 16016050 ns,
'1' after 16027000 ns, '0' after 16027050 ns,
'1' after 16038000 ns, '0' after 16038050 ns,
'1' after 16049000 ns, '0' after 16049050 ns,
'1' after 16060000 ns, '0' after 16060050 ns,
'1' after 16071000 ns, '0' after 16071050 ns,
'1' after 16082000 ns, '0' after 16082050 ns,
'1' after 16093000 ns, '0' after 16093050 ns,
'1' after 16104000 ns, '0' after 16104050 ns,
'1' after 16115000 ns, '0' after 16115050 ns,
'1' after 16126000 ns, '0' after 16126050 ns,
'1' after 16137000 ns, '0' after 16137050 ns,
'1' after 16148000 ns, '0' after 16148050 ns,
'1' after 16159000 ns, '0' after 16159050 ns,
'1' after 16170000 ns, '0' after 16170050 ns,
'1' after 16181000 ns, '0' after 16181050 ns,
'1' after 16192000 ns, '0' after 16192050 ns,
'1' after 16203000 ns, '0' after 16203050 ns,
'1' after 16214000 ns, '0' after 16214050 ns,
'1' after 16225000 ns, '0' after 16225050 ns,
'1' after 16236000 ns, '0' after 16236050 ns,
'1' after 16247000 ns, '0' after 16247050 ns,
'1' after 16258000 ns, '0' after 16258050 ns,
'1' after 16269000 ns, '0' after 16269050 ns,
'1' after 16280000 ns, '0' after 16280050 ns,
'1' after 16291000 ns, '0' after 16291050 ns,
'1' after 16302000 ns, '0' after 16302050 ns,
'1' after 16313000 ns, '0' after 16313050 ns,
'1' after 16324000 ns, '0' after 16324050 ns,
'1' after 16335000 ns, '0' after 16335050 ns,
'1' after 16346000 ns, '0' after 16346050 ns,
'1' after 16357000 ns, '0' after 16357050 ns,
'1' after 16368000 ns, '0' after 16368050 ns,
'1' after 16379000 ns, '0' after 16379050 ns,
'1' after 16390000 ns, '0' after 16390050 ns,
'1' after 16401000 ns, '0' after 16401050 ns,
'1' after 16412000 ns, '0' after 16412050 ns,
'1' after 16423000 ns, '0' after 16423050 ns,
'1' after 16434000 ns, '0' after 16434050 ns,
'1' after 16445000 ns, '0' after 16445050 ns,
'1' after 16456000 ns, '0' after 16456050 ns,
'1' after 16467000 ns, '0' after 16467050 ns,
'1' after 16478000 ns, '0' after 16478050 ns,
'1' after 16489000 ns, '0' after 16489050 ns,
'1' after 16500000 ns, '0' after 16500050 ns,
'1' after 16511000 ns, '0' after 16511050 ns,
'1' after 16522000 ns, '0' after 16522050 ns,
'1' after 16533000 ns, '0' after 16533050 ns,
'1' after 16544000 ns, '0' after 16544050 ns,
'1' after 16555000 ns, '0' after 16555050 ns,
'1' after 16566000 ns, '0' after 16566050 ns,
'1' after 16577000 ns, '0' after 16577050 ns,
'1' after 16588000 ns, '0' after 16588050 ns,
'1' after 16599000 ns, '0' after 16599050 ns,
'1' after 16610000 ns, '0' after 16610050 ns,
'1' after 16621000 ns, '0' after 16621050 ns,
'1' after 16632000 ns, '0' after 16632050 ns,
'1' after 16643000 ns, '0' after 16643050 ns,
'1' after 16654000 ns, '0' after 16654050 ns,
'1' after 16665000 ns, '0' after 16665050 ns,
'1' after 16676000 ns, '0' after 16676050 ns,
'1' after 16687000 ns, '0' after 16687050 ns,
'1' after 16698000 ns, '0' after 16698050 ns,
'1' after 16709000 ns, '0' after 16709050 ns,
'1' after 16720000 ns, '0' after 16720050 ns,
'1' after 16731000 ns, '0' after 16731050 ns,
'1' after 16742000 ns, '0' after 16742050 ns,
'1' after 16753000 ns, '0' after 16753050 ns,
'1' after 16764000 ns, '0' after 16764050 ns,
'1' after 16775000 ns, '0' after 16775050 ns,
'1' after 16786000 ns, '0' after 16786050 ns,
'1' after 16797000 ns, '0' after 16797050 ns,
'1' after 16808000 ns, '0' after 16808050 ns,
'1' after 16819000 ns, '0' after 16819050 ns,
'1' after 16830000 ns, '0' after 16830050 ns,
'1' after 16841000 ns, '0' after 16841050 ns,
'1' after 16852000 ns, '0' after 16852050 ns,
'1' after 16863000 ns, '0' after 16863050 ns,
'1' after 16874000 ns, '0' after 16874050 ns,
'1' after 16885000 ns, '0' after 16885050 ns,
'1' after 16896000 ns, '0' after 16896050 ns,
'1' after 16907000 ns, '0' after 16907050 ns,
'1' after 16918000 ns, '0' after 16918050 ns,
'1' after 16929000 ns, '0' after 16929050 ns,
'1' after 16940000 ns, '0' after 16940050 ns,
'1' after 16951000 ns, '0' after 16951050 ns,
'1' after 16962000 ns, '0' after 16962050 ns,
'1' after 16973000 ns, '0' after 16973050 ns,
'1' after 16984000 ns, '0' after 16984050 ns,
'1' after 16995000 ns, '0' after 16995050 ns,
'1' after 17006000 ns, '0' after 17006050 ns,
'1' after 17017000 ns, '0' after 17017050 ns,
'1' after 17028000 ns, '0' after 17028050 ns,
'1' after 17039000 ns, '0' after 17039050 ns,
'1' after 17050000 ns, '0' after 17050050 ns,
'1' after 17061000 ns, '0' after 17061050 ns,
'1' after 17072000 ns, '0' after 17072050 ns,
'1' after 17083000 ns, '0' after 17083050 ns,
'1' after 17094000 ns, '0' after 17094050 ns,
'1' after 17105000 ns, '0' after 17105050 ns,
'1' after 17116000 ns, '0' after 17116050 ns,
'1' after 17127000 ns, '0' after 17127050 ns,
'1' after 17138000 ns, '0' after 17138050 ns,
'1' after 17149000 ns, '0' after 17149050 ns,
'1' after 17160000 ns, '0' after 17160050 ns,
'1' after 17171000 ns, '0' after 17171050 ns,
'1' after 17182000 ns, '0' after 17182050 ns,
'1' after 17193000 ns, '0' after 17193050 ns,
'1' after 17204000 ns, '0' after 17204050 ns,
'1' after 17215000 ns, '0' after 17215050 ns,
'1' after 17226000 ns, '0' after 17226050 ns,
'1' after 17237000 ns, '0' after 17237050 ns,
'1' after 17248000 ns, '0' after 17248050 ns,
'1' after 17259000 ns, '0' after 17259050 ns,
'1' after 17270000 ns, '0' after 17270050 ns,
'1' after 17281000 ns, '0' after 17281050 ns,
'1' after 17292000 ns, '0' after 17292050 ns,
'1' after 17303000 ns, '0' after 17303050 ns,
'1' after 17314000 ns, '0' after 17314050 ns,
'1' after 17325000 ns, '0' after 17325050 ns,
'1' after 17336000 ns, '0' after 17336050 ns,
'1' after 17347000 ns, '0' after 17347050 ns,
'1' after 17358000 ns, '0' after 17358050 ns,
'1' after 17369000 ns, '0' after 17369050 ns,
'1' after 17380000 ns, '0' after 17380050 ns,
'1' after 17391000 ns, '0' after 17391050 ns,
'1' after 17402000 ns, '0' after 17402050 ns,
'1' after 17413000 ns, '0' after 17413050 ns,
'1' after 17424000 ns, '0' after 17424050 ns,
'1' after 17435000 ns, '0' after 17435050 ns,
'1' after 17446000 ns, '0' after 17446050 ns,
'1' after 17457000 ns, '0' after 17457050 ns,
'1' after 17468000 ns, '0' after 17468050 ns,
'1' after 17479000 ns, '0' after 17479050 ns,
'1' after 17490000 ns, '0' after 17490050 ns,
'1' after 17501000 ns, '0' after 17501050 ns,
'1' after 17512000 ns, '0' after 17512050 ns,
'1' after 17523000 ns, '0' after 17523050 ns,
'1' after 17534000 ns, '0' after 17534050 ns,
'1' after 17545000 ns, '0' after 17545050 ns,
'1' after 17556000 ns, '0' after 17556050 ns,
'1' after 17567000 ns, '0' after 17567050 ns,
'1' after 17578000 ns, '0' after 17578050 ns,
'1' after 17589000 ns, '0' after 17589050 ns,
'1' after 17600000 ns, '0' after 17600050 ns,
'1' after 17611000 ns, '0' after 17611050 ns,
'1' after 17622000 ns, '0' after 17622050 ns,
'1' after 17633000 ns, '0' after 17633050 ns,
'1' after 17644000 ns, '0' after 17644050 ns,
'1' after 17655000 ns, '0' after 17655050 ns,
'1' after 17666000 ns, '0' after 17666050 ns,
'1' after 17677000 ns, '0' after 17677050 ns,
'1' after 17688000 ns, '0' after 17688050 ns,
'1' after 17699000 ns, '0' after 17699050 ns,
'1' after 17710000 ns, '0' after 17710050 ns,
'1' after 17721000 ns, '0' after 17721050 ns,
'1' after 17732000 ns, '0' after 17732050 ns,
'1' after 17743000 ns, '0' after 17743050 ns,
'1' after 17754000 ns, '0' after 17754050 ns,
'1' after 17765000 ns, '0' after 17765050 ns,
'1' after 17776000 ns, '0' after 17776050 ns,
'1' after 17787000 ns, '0' after 17787050 ns,
'1' after 17798000 ns, '0' after 17798050 ns,
'1' after 17809000 ns, '0' after 17809050 ns,
'1' after 17820000 ns, '0' after 17820050 ns,
'1' after 17831000 ns, '0' after 17831050 ns,
'1' after 17842000 ns, '0' after 17842050 ns,
'1' after 17853000 ns, '0' after 17853050 ns,
'1' after 17864000 ns, '0' after 17864050 ns,
'1' after 17875000 ns, '0' after 17875050 ns,
'1' after 17886000 ns, '0' after 17886050 ns,
'1' after 17897000 ns, '0' after 17897050 ns,
'1' after 17908000 ns, '0' after 17908050 ns,
'1' after 17919000 ns, '0' after 17919050 ns,
'1' after 17930000 ns, '0' after 17930050 ns,
'1' after 17941000 ns, '0' after 17941050 ns,
'1' after 17952000 ns, '0' after 17952050 ns,
'1' after 17963000 ns, '0' after 17963050 ns,
'1' after 17974000 ns, '0' after 17974050 ns,
'1' after 17985000 ns, '0' after 17985050 ns,
'1' after 17996000 ns, '0' after 17996050 ns,
'1' after 18007000 ns, '0' after 18007050 ns,
'1' after 18018000 ns, '0' after 18018050 ns,
'1' after 18029000 ns, '0' after 18029050 ns,
'1' after 18040000 ns, '0' after 18040050 ns,
'1' after 18051000 ns, '0' after 18051050 ns,
'1' after 18062000 ns, '0' after 18062050 ns,
'1' after 18073000 ns, '0' after 18073050 ns,
'1' after 18084000 ns, '0' after 18084050 ns,
'1' after 18095000 ns, '0' after 18095050 ns,
'1' after 18106000 ns, '0' after 18106050 ns,
'1' after 18117000 ns, '0' after 18117050 ns,
'1' after 18128000 ns, '0' after 18128050 ns,
'1' after 18139000 ns, '0' after 18139050 ns,
'1' after 18150000 ns, '0' after 18150050 ns,
'1' after 18161000 ns, '0' after 18161050 ns,
'1' after 18172000 ns, '0' after 18172050 ns,
'1' after 18183000 ns, '0' after 18183050 ns,
'1' after 18194000 ns, '0' after 18194050 ns,
'1' after 18205000 ns, '0' after 18205050 ns,
'1' after 18216000 ns, '0' after 18216050 ns,
'1' after 18227000 ns, '0' after 18227050 ns,
'1' after 18238000 ns, '0' after 18238050 ns,
'1' after 18249000 ns, '0' after 18249050 ns,
'1' after 18260000 ns, '0' after 18260050 ns,
'1' after 18271000 ns, '0' after 18271050 ns,
'1' after 18282000 ns, '0' after 18282050 ns,
'1' after 18293000 ns, '0' after 18293050 ns,
'1' after 18304000 ns, '0' after 18304050 ns,
'1' after 18315000 ns, '0' after 18315050 ns,
'1' after 18326000 ns, '0' after 18326050 ns,
'1' after 18337000 ns, '0' after 18337050 ns,
'1' after 18348000 ns, '0' after 18348050 ns,
'1' after 18359000 ns, '0' after 18359050 ns,
'1' after 18370000 ns, '0' after 18370050 ns,
'1' after 18381000 ns, '0' after 18381050 ns,
'1' after 18392000 ns, '0' after 18392050 ns,
'1' after 18403000 ns, '0' after 18403050 ns,
'1' after 18414000 ns, '0' after 18414050 ns,
'1' after 18425000 ns, '0' after 18425050 ns,
'1' after 18436000 ns, '0' after 18436050 ns,
'1' after 18447000 ns, '0' after 18447050 ns,
'1' after 18458000 ns, '0' after 18458050 ns,
'1' after 18469000 ns, '0' after 18469050 ns,
'1' after 18480000 ns, '0' after 18480050 ns,
'1' after 18491000 ns, '0' after 18491050 ns,
'1' after 18502000 ns, '0' after 18502050 ns,
'1' after 18513000 ns, '0' after 18513050 ns,
'1' after 18524000 ns, '0' after 18524050 ns,
'1' after 18535000 ns, '0' after 18535050 ns,
'1' after 18546000 ns, '0' after 18546050 ns,
'1' after 18557000 ns, '0' after 18557050 ns,
'1' after 18568000 ns, '0' after 18568050 ns,
'1' after 18579000 ns, '0' after 18579050 ns,
'1' after 18590000 ns, '0' after 18590050 ns,
'1' after 18601000 ns, '0' after 18601050 ns,
'1' after 18612000 ns, '0' after 18612050 ns,
'1' after 18623000 ns, '0' after 18623050 ns,
'1' after 18634000 ns, '0' after 18634050 ns,
'1' after 18645000 ns, '0' after 18645050 ns,
'1' after 18656000 ns, '0' after 18656050 ns,
'1' after 18667000 ns, '0' after 18667050 ns,
'1' after 18678000 ns, '0' after 18678050 ns,
'1' after 18689000 ns, '0' after 18689050 ns,
'1' after 18700000 ns, '0' after 18700050 ns,
'1' after 18711000 ns, '0' after 18711050 ns,
'1' after 18722000 ns, '0' after 18722050 ns,
'1' after 18733000 ns, '0' after 18733050 ns,
'1' after 18744000 ns, '0' after 18744050 ns,
'1' after 18755000 ns, '0' after 18755050 ns,
'1' after 18766000 ns, '0' after 18766050 ns,
'1' after 18777000 ns, '0' after 18777050 ns,
'1' after 18788000 ns, '0' after 18788050 ns,
'1' after 18799000 ns, '0' after 18799050 ns,
'1' after 18810000 ns, '0' after 18810050 ns,
'1' after 18821000 ns, '0' after 18821050 ns,
'1' after 18832000 ns, '0' after 18832050 ns,
'1' after 18843000 ns, '0' after 18843050 ns,
'1' after 18854000 ns, '0' after 18854050 ns,
'1' after 18865000 ns, '0' after 18865050 ns,
'1' after 18876000 ns, '0' after 18876050 ns,
'1' after 18887000 ns, '0' after 18887050 ns,
'1' after 18898000 ns, '0' after 18898050 ns,
'1' after 18909000 ns, '0' after 18909050 ns,
'1' after 18920000 ns, '0' after 18920050 ns,
'1' after 18931000 ns, '0' after 18931050 ns,
'1' after 18942000 ns, '0' after 18942050 ns,
'1' after 18953000 ns, '0' after 18953050 ns,
'1' after 18964000 ns, '0' after 18964050 ns,
'1' after 18975000 ns, '0' after 18975050 ns,
'1' after 18986000 ns, '0' after 18986050 ns,
'1' after 18997000 ns, '0' after 18997050 ns,
'1' after 19008000 ns, '0' after 19008050 ns,
'1' after 19019000 ns, '0' after 19019050 ns,
'1' after 19030000 ns, '0' after 19030050 ns,
'1' after 19041000 ns, '0' after 19041050 ns,
'1' after 19052000 ns, '0' after 19052050 ns,
'1' after 19063000 ns, '0' after 19063050 ns,
'1' after 19074000 ns, '0' after 19074050 ns,
'1' after 19085000 ns, '0' after 19085050 ns,
'1' after 19096000 ns, '0' after 19096050 ns,
'1' after 19107000 ns, '0' after 19107050 ns,
'1' after 19118000 ns, '0' after 19118050 ns,
'1' after 19129000 ns, '0' after 19129050 ns,
'1' after 19140000 ns, '0' after 19140050 ns,
'1' after 19151000 ns, '0' after 19151050 ns,
'1' after 19162000 ns, '0' after 19162050 ns,
'1' after 19173000 ns, '0' after 19173050 ns,
'1' after 19184000 ns, '0' after 19184050 ns,
'1' after 19195000 ns, '0' after 19195050 ns,
'1' after 19206000 ns, '0' after 19206050 ns,
'1' after 19217000 ns, '0' after 19217050 ns,
'1' after 19228000 ns, '0' after 19228050 ns,
'1' after 19239000 ns, '0' after 19239050 ns,
'1' after 19250000 ns, '0' after 19250050 ns,
'1' after 19261000 ns, '0' after 19261050 ns,
'1' after 19272000 ns, '0' after 19272050 ns,
'1' after 19283000 ns, '0' after 19283050 ns,
'1' after 19294000 ns, '0' after 19294050 ns,
'1' after 19305000 ns, '0' after 19305050 ns,
'1' after 19316000 ns, '0' after 19316050 ns,
'1' after 19327000 ns, '0' after 19327050 ns,
'1' after 19338000 ns, '0' after 19338050 ns,
'1' after 19349000 ns, '0' after 19349050 ns,
'1' after 19360000 ns, '0' after 19360050 ns,
'1' after 19371000 ns, '0' after 19371050 ns,
'1' after 19382000 ns, '0' after 19382050 ns,
'1' after 19393000 ns, '0' after 19393050 ns,
'1' after 19404000 ns, '0' after 19404050 ns,
'1' after 19415000 ns, '0' after 19415050 ns,
'1' after 19426000 ns, '0' after 19426050 ns,
'1' after 19437000 ns, '0' after 19437050 ns,
'1' after 19448000 ns, '0' after 19448050 ns,
'1' after 19459000 ns, '0' after 19459050 ns,
'1' after 19470000 ns, '0' after 19470050 ns,
'1' after 19481000 ns, '0' after 19481050 ns,
'1' after 19492000 ns, '0' after 19492050 ns,
'1' after 19503000 ns, '0' after 19503050 ns,
'1' after 19514000 ns, '0' after 19514050 ns,
'1' after 19525000 ns, '0' after 19525050 ns,
'1' after 19536000 ns, '0' after 19536050 ns,
'1' after 19547000 ns, '0' after 19547050 ns,
'1' after 19558000 ns, '0' after 19558050 ns,
'1' after 19569000 ns, '0' after 19569050 ns,
'1' after 19580000 ns, '0' after 19580050 ns,
'1' after 19591000 ns, '0' after 19591050 ns,
'1' after 19602000 ns, '0' after 19602050 ns,
'1' after 19613000 ns, '0' after 19613050 ns,
'1' after 19624000 ns, '0' after 19624050 ns,
'1' after 19635000 ns, '0' after 19635050 ns,
'1' after 19646000 ns, '0' after 19646050 ns,
'1' after 19657000 ns, '0' after 19657050 ns,
'1' after 19668000 ns, '0' after 19668050 ns,
'1' after 19679000 ns, '0' after 19679050 ns,
'1' after 19690000 ns, '0' after 19690050 ns,
'1' after 19701000 ns, '0' after 19701050 ns,
'1' after 19712000 ns, '0' after 19712050 ns,
'1' after 19723000 ns, '0' after 19723050 ns,
'1' after 19734000 ns, '0' after 19734050 ns,
'1' after 19745000 ns, '0' after 19745050 ns,
'1' after 19756000 ns, '0' after 19756050 ns,
'1' after 19767000 ns, '0' after 19767050 ns,
'1' after 19778000 ns, '0' after 19778050 ns,
'1' after 19789000 ns, '0' after 19789050 ns,
'1' after 19800000 ns, '0' after 19800050 ns,
'1' after 19811000 ns, '0' after 19811050 ns,
'1' after 19822000 ns, '0' after 19822050 ns,
'1' after 19833000 ns, '0' after 19833050 ns,
'1' after 19844000 ns, '0' after 19844050 ns,
'1' after 19855000 ns, '0' after 19855050 ns,
'1' after 19866000 ns, '0' after 19866050 ns,
'1' after 19877000 ns, '0' after 19877050 ns,
'1' after 19888000 ns, '0' after 19888050 ns,
'1' after 19899000 ns, '0' after 19899050 ns,
'1' after 19910000 ns, '0' after 19910050 ns,
'1' after 19921000 ns, '0' after 19921050 ns,
'1' after 19932000 ns, '0' after 19932050 ns,
'1' after 19943000 ns, '0' after 19943050 ns,
'1' after 19954000 ns, '0' after 19954050 ns,
'1' after 19965000 ns, '0' after 19965050 ns,
'1' after 19976000 ns, '0' after 19976050 ns,
'1' after 19987000 ns, '0' after 19987050 ns,
'1' after 19998000 ns, '0' after 19998050 ns,
'1' after 20009000 ns, '0' after 20009050 ns,
'1' after 20020000 ns, '0' after 20020050 ns,
'1' after 20031000 ns, '0' after 20031050 ns,
'1' after 20042000 ns, '0' after 20042050 ns,
'1' after 20053000 ns, '0' after 20053050 ns,
'1' after 20064000 ns, '0' after 20064050 ns,
'1' after 20075000 ns, '0' after 20075050 ns,
'1' after 20086000 ns, '0' after 20086050 ns,
'1' after 20097000 ns, '0' after 20097050 ns,
'1' after 20108000 ns, '0' after 20108050 ns,
'1' after 20119000 ns, '0' after 20119050 ns,
'1' after 20130000 ns, '0' after 20130050 ns,
'1' after 20141000 ns, '0' after 20141050 ns,
'1' after 20152000 ns, '0' after 20152050 ns,
'1' after 20163000 ns, '0' after 20163050 ns,
'1' after 20174000 ns, '0' after 20174050 ns,
'1' after 20185000 ns, '0' after 20185050 ns,
'1' after 20196000 ns, '0' after 20196050 ns,
'1' after 20207000 ns, '0' after 20207050 ns,
'1' after 20218000 ns, '0' after 20218050 ns,
'1' after 20229000 ns, '0' after 20229050 ns,
'1' after 20240000 ns, '0' after 20240050 ns,
'1' after 20251000 ns, '0' after 20251050 ns,
'1' after 20262000 ns, '0' after 20262050 ns,
'1' after 20273000 ns, '0' after 20273050 ns,
'1' after 20284000 ns, '0' after 20284050 ns,
'1' after 20295000 ns, '0' after 20295050 ns,
'1' after 20306000 ns, '0' after 20306050 ns,
'1' after 20317000 ns, '0' after 20317050 ns,
'1' after 20328000 ns, '0' after 20328050 ns,
'1' after 20339000 ns, '0' after 20339050 ns,
'1' after 20350000 ns, '0' after 20350050 ns,
'1' after 20361000 ns, '0' after 20361050 ns,
'1' after 20372000 ns, '0' after 20372050 ns,
'1' after 20383000 ns, '0' after 20383050 ns,
'1' after 20394000 ns, '0' after 20394050 ns,
'1' after 20405000 ns, '0' after 20405050 ns,
'1' after 20416000 ns, '0' after 20416050 ns,
'1' after 20427000 ns, '0' after 20427050 ns,
'1' after 20438000 ns, '0' after 20438050 ns,
'1' after 20449000 ns, '0' after 20449050 ns,
'1' after 20460000 ns, '0' after 20460050 ns,
'1' after 20471000 ns, '0' after 20471050 ns,
'1' after 20482000 ns, '0' after 20482050 ns,
'1' after 20493000 ns, '0' after 20493050 ns,
'1' after 20504000 ns, '0' after 20504050 ns,
'1' after 20515000 ns, '0' after 20515050 ns,
'1' after 20526000 ns, '0' after 20526050 ns,
'1' after 20537000 ns, '0' after 20537050 ns,
'1' after 20548000 ns, '0' after 20548050 ns,
'1' after 20559000 ns, '0' after 20559050 ns,
'1' after 20570000 ns, '0' after 20570050 ns,
'1' after 20581000 ns, '0' after 20581050 ns,
'1' after 20592000 ns, '0' after 20592050 ns,
'1' after 20603000 ns, '0' after 20603050 ns,
'1' after 20614000 ns, '0' after 20614050 ns,
'1' after 20625000 ns, '0' after 20625050 ns,
'1' after 20636000 ns, '0' after 20636050 ns,
'1' after 20647000 ns, '0' after 20647050 ns,
'1' after 20658000 ns, '0' after 20658050 ns,
'1' after 20669000 ns, '0' after 20669050 ns,
'1' after 20680000 ns, '0' after 20680050 ns,
'1' after 20691000 ns, '0' after 20691050 ns,
'1' after 20702000 ns, '0' after 20702050 ns,
'1' after 20713000 ns, '0' after 20713050 ns,
'1' after 20724000 ns, '0' after 20724050 ns,
'1' after 20735000 ns, '0' after 20735050 ns,
'1' after 20746000 ns, '0' after 20746050 ns,
'1' after 20757000 ns, '0' after 20757050 ns,
'1' after 20768000 ns, '0' after 20768050 ns,
'1' after 20779000 ns, '0' after 20779050 ns,
'1' after 20790000 ns, '0' after 20790050 ns,
'1' after 20801000 ns, '0' after 20801050 ns,
'1' after 20812000 ns, '0' after 20812050 ns,
'1' after 20823000 ns, '0' after 20823050 ns,
'1' after 20834000 ns, '0' after 20834050 ns,
'1' after 20845000 ns, '0' after 20845050 ns,
'1' after 20856000 ns, '0' after 20856050 ns,
'1' after 20867000 ns, '0' after 20867050 ns,
'1' after 20878000 ns, '0' after 20878050 ns,
'1' after 20889000 ns, '0' after 20889050 ns,
'1' after 20900000 ns, '0' after 20900050 ns,
'1' after 20911000 ns, '0' after 20911050 ns,
'1' after 20922000 ns, '0' after 20922050 ns,
'1' after 20933000 ns, '0' after 20933050 ns,
'1' after 20944000 ns, '0' after 20944050 ns,
'1' after 20955000 ns, '0' after 20955050 ns,
'1' after 20966000 ns, '0' after 20966050 ns,
'1' after 20977000 ns, '0' after 20977050 ns,
'1' after 20988000 ns, '0' after 20988050 ns,
'1' after 20999000 ns, '0' after 20999050 ns,
'1' after 21010000 ns, '0' after 21010050 ns,
'1' after 21021000 ns, '0' after 21021050 ns,
'1' after 21032000 ns, '0' after 21032050 ns,
'1' after 21043000 ns, '0' after 21043050 ns,
'1' after 21054000 ns, '0' after 21054050 ns,
'1' after 21065000 ns, '0' after 21065050 ns,
'1' after 21076000 ns, '0' after 21076050 ns,
'1' after 21087000 ns, '0' after 21087050 ns,
'1' after 21098000 ns, '0' after 21098050 ns,
'1' after 21109000 ns, '0' after 21109050 ns,
'1' after 21120000 ns, '0' after 21120050 ns,
'1' after 21131000 ns, '0' after 21131050 ns,
'1' after 21142000 ns, '0' after 21142050 ns,
'1' after 21153000 ns, '0' after 21153050 ns,
'1' after 21164000 ns, '0' after 21164050 ns,
'1' after 21175000 ns, '0' after 21175050 ns,
'1' after 21186000 ns, '0' after 21186050 ns,
'1' after 21197000 ns, '0' after 21197050 ns,
'1' after 21208000 ns, '0' after 21208050 ns,
'1' after 21219000 ns, '0' after 21219050 ns,
'1' after 21230000 ns, '0' after 21230050 ns,
'1' after 21241000 ns, '0' after 21241050 ns,
'1' after 21252000 ns, '0' after 21252050 ns,
'1' after 21263000 ns, '0' after 21263050 ns,
'1' after 21274000 ns, '0' after 21274050 ns,
'1' after 21285000 ns, '0' after 21285050 ns,
'1' after 21296000 ns, '0' after 21296050 ns,
'1' after 21307000 ns, '0' after 21307050 ns,
'1' after 21318000 ns, '0' after 21318050 ns,
'1' after 21329000 ns, '0' after 21329050 ns,
'1' after 21340000 ns, '0' after 21340050 ns,
'1' after 21351000 ns, '0' after 21351050 ns,
'1' after 21362000 ns, '0' after 21362050 ns,
'1' after 21373000 ns, '0' after 21373050 ns,
'1' after 21384000 ns, '0' after 21384050 ns,
'1' after 21395000 ns, '0' after 21395050 ns,
'1' after 21406000 ns, '0' after 21406050 ns,
'1' after 21417000 ns, '0' after 21417050 ns,
'1' after 21428000 ns, '0' after 21428050 ns,
'1' after 21439000 ns, '0' after 21439050 ns,
'1' after 21450000 ns, '0' after 21450050 ns,
'1' after 21461000 ns, '0' after 21461050 ns,
'1' after 21472000 ns, '0' after 21472050 ns,
'1' after 21483000 ns, '0' after 21483050 ns,
'1' after 21494000 ns, '0' after 21494050 ns,
'1' after 21505000 ns, '0' after 21505050 ns,
'1' after 21516000 ns, '0' after 21516050 ns,
'1' after 21527000 ns, '0' after 21527050 ns,
'1' after 21538000 ns, '0' after 21538050 ns,
'1' after 21549000 ns, '0' after 21549050 ns,
'1' after 21560000 ns, '0' after 21560050 ns,
'1' after 21571000 ns, '0' after 21571050 ns,
'1' after 21582000 ns, '0' after 21582050 ns,
'1' after 21593000 ns, '0' after 21593050 ns,
'1' after 21604000 ns, '0' after 21604050 ns,
'1' after 21615000 ns, '0' after 21615050 ns,
'1' after 21626000 ns, '0' after 21626050 ns,
'1' after 21637000 ns, '0' after 21637050 ns,
'1' after 21648000 ns, '0' after 21648050 ns,
'1' after 21659000 ns, '0' after 21659050 ns,
'1' after 21670000 ns, '0' after 21670050 ns,
'1' after 21681000 ns, '0' after 21681050 ns,
'1' after 21692000 ns, '0' after 21692050 ns,
'1' after 21703000 ns, '0' after 21703050 ns,
'1' after 21714000 ns, '0' after 21714050 ns,
'1' after 21725000 ns, '0' after 21725050 ns,
'1' after 21736000 ns, '0' after 21736050 ns,
'1' after 21747000 ns, '0' after 21747050 ns,
'1' after 21758000 ns, '0' after 21758050 ns,
'1' after 21769000 ns, '0' after 21769050 ns,
'1' after 21780000 ns, '0' after 21780050 ns,
'1' after 21791000 ns, '0' after 21791050 ns,
'1' after 21802000 ns, '0' after 21802050 ns,
'1' after 21813000 ns, '0' after 21813050 ns,
'1' after 21824000 ns, '0' after 21824050 ns,
'1' after 21835000 ns, '0' after 21835050 ns,
'1' after 21846000 ns, '0' after 21846050 ns,
'1' after 21857000 ns, '0' after 21857050 ns,
'1' after 21868000 ns, '0' after 21868050 ns,
'1' after 21879000 ns, '0' after 21879050 ns,
'1' after 21890000 ns, '0' after 21890050 ns,
'1' after 21901000 ns, '0' after 21901050 ns,
'1' after 21912000 ns, '0' after 21912050 ns,
'1' after 21923000 ns, '0' after 21923050 ns,
'1' after 21934000 ns, '0' after 21934050 ns,
'1' after 21945000 ns, '0' after 21945050 ns,
'1' after 21956000 ns, '0' after 21956050 ns,
'1' after 21967000 ns, '0' after 21967050 ns,
'1' after 21978000 ns, '0' after 21978050 ns,
'1' after 21989000 ns, '0' after 21989050 ns,
'1' after 22000000 ns, '0' after 22000050 ns,
'1' after 22011000 ns, '0' after 22011050 ns,
'1' after 22022000 ns, '0' after 22022050 ns,
'1' after 22033000 ns, '0' after 22033050 ns,
'1' after 22044000 ns, '0' after 22044050 ns,
'1' after 22055000 ns, '0' after 22055050 ns,
'1' after 22066000 ns, '0' after 22066050 ns,
'1' after 22077000 ns, '0' after 22077050 ns,
'1' after 22088000 ns, '0' after 22088050 ns,
'1' after 22099000 ns, '0' after 22099050 ns,
'1' after 22110000 ns, '0' after 22110050 ns,
'1' after 22121000 ns, '0' after 22121050 ns,
'1' after 22132000 ns, '0' after 22132050 ns,
'1' after 22143000 ns, '0' after 22143050 ns,
'1' after 22154000 ns, '0' after 22154050 ns,
'1' after 22165000 ns, '0' after 22165050 ns,
'1' after 22176000 ns, '0' after 22176050 ns,
'1' after 22187000 ns, '0' after 22187050 ns,
'1' after 22198000 ns, '0' after 22198050 ns,
'1' after 22209000 ns, '0' after 22209050 ns,
'1' after 22220000 ns, '0' after 22220050 ns,
'1' after 22231000 ns, '0' after 22231050 ns,
'1' after 22242000 ns, '0' after 22242050 ns,
'1' after 22253000 ns, '0' after 22253050 ns,
'1' after 22264000 ns, '0' after 22264050 ns,
'1' after 22275000 ns, '0' after 22275050 ns,
'1' after 22286000 ns, '0' after 22286050 ns,
'1' after 22297000 ns, '0' after 22297050 ns,
'1' after 22308000 ns, '0' after 22308050 ns,
'1' after 22319000 ns, '0' after 22319050 ns,
'1' after 22330000 ns, '0' after 22330050 ns,
'1' after 22341000 ns, '0' after 22341050 ns,
'1' after 22352000 ns, '0' after 22352050 ns,
'1' after 22363000 ns, '0' after 22363050 ns,
'1' after 22374000 ns, '0' after 22374050 ns,
'1' after 22385000 ns, '0' after 22385050 ns,
'1' after 22396000 ns, '0' after 22396050 ns,
'1' after 22407000 ns, '0' after 22407050 ns,
'1' after 22418000 ns, '0' after 22418050 ns,
'1' after 22429000 ns, '0' after 22429050 ns,
'1' after 22440000 ns, '0' after 22440050 ns,
'1' after 22451000 ns, '0' after 22451050 ns,
'1' after 22462000 ns, '0' after 22462050 ns,
'1' after 22473000 ns, '0' after 22473050 ns,
'1' after 22484000 ns, '0' after 22484050 ns,
'1' after 22495000 ns, '0' after 22495050 ns,
'1' after 22506000 ns, '0' after 22506050 ns,
'1' after 22517000 ns, '0' after 22517050 ns,
'1' after 22528000 ns, '0' after 22528050 ns,
'1' after 22539000 ns, '0' after 22539050 ns,
'1' after 22550000 ns, '0' after 22550050 ns,
'1' after 22561000 ns, '0' after 22561050 ns,
'1' after 22572000 ns, '0' after 22572050 ns,
'1' after 22583000 ns, '0' after 22583050 ns,
'1' after 22594000 ns, '0' after 22594050 ns,
'1' after 22605000 ns, '0' after 22605050 ns,
'1' after 22616000 ns, '0' after 22616050 ns,
'1' after 22627000 ns, '0' after 22627050 ns,
'1' after 22638000 ns, '0' after 22638050 ns,
'1' after 22649000 ns, '0' after 22649050 ns,
'1' after 22660000 ns, '0' after 22660050 ns,
'1' after 22671000 ns, '0' after 22671050 ns,
'1' after 22682000 ns, '0' after 22682050 ns,
'1' after 22693000 ns, '0' after 22693050 ns,
'1' after 22704000 ns, '0' after 22704050 ns,
'1' after 22715000 ns, '0' after 22715050 ns,
'1' after 22726000 ns, '0' after 22726050 ns,
'1' after 22737000 ns, '0' after 22737050 ns,
'1' after 22748000 ns, '0' after 22748050 ns,
'1' after 22759000 ns, '0' after 22759050 ns,
'1' after 22770000 ns, '0' after 22770050 ns,
'1' after 22781000 ns, '0' after 22781050 ns,
'1' after 22792000 ns, '0' after 22792050 ns,
'1' after 22803000 ns, '0' after 22803050 ns,
'1' after 22814000 ns, '0' after 22814050 ns,
'1' after 22825000 ns, '0' after 22825050 ns,
'1' after 22836000 ns, '0' after 22836050 ns,
'1' after 22847000 ns, '0' after 22847050 ns,
'1' after 22858000 ns, '0' after 22858050 ns,
'1' after 22869000 ns, '0' after 22869050 ns,
'1' after 22880000 ns, '0' after 22880050 ns,
'1' after 22891000 ns, '0' after 22891050 ns,
'1' after 22902000 ns, '0' after 22902050 ns,
'1' after 22913000 ns, '0' after 22913050 ns,
'1' after 22924000 ns, '0' after 22924050 ns,
'1' after 22935000 ns, '0' after 22935050 ns,
'1' after 22946000 ns, '0' after 22946050 ns,
'1' after 22957000 ns, '0' after 22957050 ns,
'1' after 22968000 ns, '0' after 22968050 ns,
'1' after 22979000 ns, '0' after 22979050 ns,
'1' after 22990000 ns, '0' after 22990050 ns,
'1' after 23001000 ns, '0' after 23001050 ns,
'1' after 23012000 ns, '0' after 23012050 ns,
'1' after 23023000 ns, '0' after 23023050 ns,
'1' after 23034000 ns, '0' after 23034050 ns,
'1' after 23045000 ns, '0' after 23045050 ns,
'1' after 23056000 ns, '0' after 23056050 ns,
'1' after 23067000 ns, '0' after 23067050 ns,
'1' after 23078000 ns, '0' after 23078050 ns,
'1' after 23089000 ns, '0' after 23089050 ns,
'1' after 23100000 ns, '0' after 23100050 ns,
'1' after 23111000 ns, '0' after 23111050 ns,
'1' after 23122000 ns, '0' after 23122050 ns,
'1' after 23133000 ns, '0' after 23133050 ns,
'1' after 23144000 ns, '0' after 23144050 ns,
'1' after 23155000 ns, '0' after 23155050 ns,
'1' after 23166000 ns, '0' after 23166050 ns,
'1' after 23177000 ns, '0' after 23177050 ns,
'1' after 23188000 ns, '0' after 23188050 ns,
'1' after 23199000 ns, '0' after 23199050 ns,
'1' after 23210000 ns, '0' after 23210050 ns,
'1' after 23221000 ns, '0' after 23221050 ns,
'1' after 23232000 ns, '0' after 23232050 ns,
'1' after 23243000 ns, '0' after 23243050 ns,
'1' after 23254000 ns, '0' after 23254050 ns,
'1' after 23265000 ns, '0' after 23265050 ns,
'1' after 23276000 ns, '0' after 23276050 ns,
'1' after 23287000 ns, '0' after 23287050 ns,
'1' after 23298000 ns, '0' after 23298050 ns,
'1' after 23309000 ns, '0' after 23309050 ns,
'1' after 23320000 ns, '0' after 23320050 ns,
'1' after 23331000 ns, '0' after 23331050 ns,
'1' after 23342000 ns, '0' after 23342050 ns,
'1' after 23353000 ns, '0' after 23353050 ns,
'1' after 23364000 ns, '0' after 23364050 ns,
'1' after 23375000 ns, '0' after 23375050 ns,
'1' after 23386000 ns, '0' after 23386050 ns,
'1' after 23397000 ns, '0' after 23397050 ns,
'1' after 23408000 ns, '0' after 23408050 ns,
'1' after 23419000 ns, '0' after 23419050 ns,
'1' after 23430000 ns, '0' after 23430050 ns,
'1' after 23441000 ns, '0' after 23441050 ns,
'1' after 23452000 ns, '0' after 23452050 ns,
'1' after 23463000 ns, '0' after 23463050 ns,
'1' after 23474000 ns, '0' after 23474050 ns,
'1' after 23485000 ns, '0' after 23485050 ns,
'1' after 23496000 ns, '0' after 23496050 ns,
'1' after 23507000 ns, '0' after 23507050 ns,
'1' after 23518000 ns, '0' after 23518050 ns,
'1' after 23529000 ns, '0' after 23529050 ns,
'1' after 23540000 ns, '0' after 23540050 ns,
'1' after 23551000 ns, '0' after 23551050 ns,
'1' after 23562000 ns, '0' after 23562050 ns,
'1' after 23573000 ns, '0' after 23573050 ns,
'1' after 23584000 ns, '0' after 23584050 ns,
'1' after 23595000 ns, '0' after 23595050 ns,
'1' after 23606000 ns, '0' after 23606050 ns,
'1' after 23617000 ns, '0' after 23617050 ns,
'1' after 23628000 ns, '0' after 23628050 ns,
'1' after 23639000 ns, '0' after 23639050 ns,
'1' after 23650000 ns, '0' after 23650050 ns,
'1' after 23661000 ns, '0' after 23661050 ns,
'1' after 23672000 ns, '0' after 23672050 ns,
'1' after 23683000 ns, '0' after 23683050 ns,
'1' after 23694000 ns, '0' after 23694050 ns,
'1' after 23705000 ns, '0' after 23705050 ns,
'1' after 23716000 ns, '0' after 23716050 ns,
'1' after 23727000 ns, '0' after 23727050 ns,
'1' after 23738000 ns, '0' after 23738050 ns,
'1' after 23749000 ns, '0' after 23749050 ns,
'1' after 23760000 ns, '0' after 23760050 ns,
'1' after 23771000 ns, '0' after 23771050 ns,
'1' after 23782000 ns, '0' after 23782050 ns,
'1' after 23793000 ns, '0' after 23793050 ns,
'1' after 23804000 ns, '0' after 23804050 ns,
'1' after 23815000 ns, '0' after 23815050 ns,
'1' after 23826000 ns, '0' after 23826050 ns,
'1' after 23837000 ns, '0' after 23837050 ns,
'1' after 23848000 ns, '0' after 23848050 ns,
'1' after 23859000 ns, '0' after 23859050 ns,
'1' after 23870000 ns, '0' after 23870050 ns,
'1' after 23881000 ns, '0' after 23881050 ns,
'1' after 23892000 ns, '0' after 23892050 ns,
'1' after 23903000 ns, '0' after 23903050 ns,
'1' after 23914000 ns, '0' after 23914050 ns,
'1' after 23925000 ns, '0' after 23925050 ns,
'1' after 23936000 ns, '0' after 23936050 ns,
'1' after 23947000 ns, '0' after 23947050 ns,
'1' after 23958000 ns, '0' after 23958050 ns,
'1' after 23969000 ns, '0' after 23969050 ns,
'1' after 23980000 ns, '0' after 23980050 ns,
'1' after 23991000 ns, '0' after 23991050 ns,
'1' after 24002000 ns, '0' after 24002050 ns,
'1' after 24013000 ns, '0' after 24013050 ns,
'1' after 24024000 ns, '0' after 24024050 ns,
'1' after 24035000 ns, '0' after 24035050 ns,
'1' after 24046000 ns, '0' after 24046050 ns,
'1' after 24057000 ns, '0' after 24057050 ns,
'1' after 24068000 ns, '0' after 24068050 ns,
'1' after 24079000 ns, '0' after 24079050 ns,
'1' after 24090000 ns, '0' after 24090050 ns,
'1' after 24101000 ns, '0' after 24101050 ns,
'1' after 24112000 ns, '0' after 24112050 ns,
'1' after 24123000 ns, '0' after 24123050 ns,
'1' after 24134000 ns, '0' after 24134050 ns,
'1' after 24145000 ns, '0' after 24145050 ns,
'1' after 24156000 ns, '0' after 24156050 ns,
'1' after 24167000 ns, '0' after 24167050 ns,
'1' after 24178000 ns, '0' after 24178050 ns,
'1' after 24189000 ns, '0' after 24189050 ns,
'1' after 24200000 ns, '0' after 24200050 ns,
'1' after 24211000 ns, '0' after 24211050 ns,
'1' after 24222000 ns, '0' after 24222050 ns,
'1' after 24233000 ns, '0' after 24233050 ns,
'1' after 24244000 ns, '0' after 24244050 ns,
'1' after 24255000 ns, '0' after 24255050 ns,
'1' after 24266000 ns, '0' after 24266050 ns,
'1' after 24277000 ns, '0' after 24277050 ns,
'1' after 24288000 ns, '0' after 24288050 ns,
'1' after 24299000 ns, '0' after 24299050 ns,
'1' after 24310000 ns, '0' after 24310050 ns,
'1' after 24321000 ns, '0' after 24321050 ns,
'1' after 24332000 ns, '0' after 24332050 ns,
'1' after 24343000 ns, '0' after 24343050 ns,
'1' after 24354000 ns, '0' after 24354050 ns,
'1' after 24365000 ns, '0' after 24365050 ns,
'1' after 24376000 ns, '0' after 24376050 ns,
'1' after 24387000 ns, '0' after 24387050 ns,
'1' after 24398000 ns, '0' after 24398050 ns,
'1' after 24409000 ns, '0' after 24409050 ns,
'1' after 24420000 ns, '0' after 24420050 ns,
'1' after 24431000 ns, '0' after 24431050 ns,
'1' after 24442000 ns, '0' after 24442050 ns,
'1' after 24453000 ns, '0' after 24453050 ns,
'1' after 24464000 ns, '0' after 24464050 ns,
'1' after 24475000 ns, '0' after 24475050 ns,
'1' after 24486000 ns, '0' after 24486050 ns,
'1' after 24497000 ns, '0' after 24497050 ns,
'1' after 24508000 ns, '0' after 24508050 ns,
'1' after 24519000 ns, '0' after 24519050 ns,
'1' after 24530000 ns, '0' after 24530050 ns,
'1' after 24541000 ns, '0' after 24541050 ns,
'1' after 24552000 ns, '0' after 24552050 ns,
'1' after 24563000 ns, '0' after 24563050 ns,
'1' after 24574000 ns, '0' after 24574050 ns,
'1' after 24585000 ns, '0' after 24585050 ns,
'1' after 24596000 ns, '0' after 24596050 ns,
'1' after 24607000 ns, '0' after 24607050 ns,
'1' after 24618000 ns, '0' after 24618050 ns,
'1' after 24629000 ns, '0' after 24629050 ns,
'1' after 24640000 ns, '0' after 24640050 ns,
'1' after 24651000 ns, '0' after 24651050 ns,
'1' after 24662000 ns, '0' after 24662050 ns,
'1' after 24673000 ns, '0' after 24673050 ns,
'1' after 24684000 ns, '0' after 24684050 ns,
'1' after 24695000 ns, '0' after 24695050 ns,
'1' after 24706000 ns, '0' after 24706050 ns,
'1' after 24717000 ns, '0' after 24717050 ns,
'1' after 24728000 ns, '0' after 24728050 ns,
'1' after 24739000 ns, '0' after 24739050 ns,
'1' after 24750000 ns, '0' after 24750050 ns,
'1' after 24761000 ns, '0' after 24761050 ns,
'1' after 24772000 ns, '0' after 24772050 ns,
'1' after 24783000 ns, '0' after 24783050 ns,
'1' after 24794000 ns, '0' after 24794050 ns,
'1' after 24805000 ns, '0' after 24805050 ns,
'1' after 24816000 ns, '0' after 24816050 ns,
'1' after 24827000 ns, '0' after 24827050 ns,
'1' after 24838000 ns, '0' after 24838050 ns,
'1' after 24849000 ns, '0' after 24849050 ns,
'1' after 24860000 ns, '0' after 24860050 ns,
'1' after 24871000 ns, '0' after 24871050 ns,
'1' after 24882000 ns, '0' after 24882050 ns,
'1' after 24893000 ns, '0' after 24893050 ns,
'1' after 24904000 ns, '0' after 24904050 ns,
'1' after 24915000 ns, '0' after 24915050 ns,
'1' after 24926000 ns, '0' after 24926050 ns,
'1' after 24937000 ns, '0' after 24937050 ns,
'1' after 24948000 ns, '0' after 24948050 ns,
'1' after 24959000 ns, '0' after 24959050 ns,
'1' after 24970000 ns, '0' after 24970050 ns,
'1' after 24981000 ns, '0' after 24981050 ns,
'1' after 24992000 ns, '0' after 24992050 ns,
'1' after 25003000 ns, '0' after 25003050 ns,
'1' after 25014000 ns, '0' after 25014050 ns,
'1' after 25025000 ns, '0' after 25025050 ns,
'1' after 25036000 ns, '0' after 25036050 ns,
'1' after 25047000 ns, '0' after 25047050 ns,
'1' after 25058000 ns, '0' after 25058050 ns,
'1' after 25069000 ns, '0' after 25069050 ns,
'1' after 25080000 ns, '0' after 25080050 ns,
'1' after 25091000 ns, '0' after 25091050 ns,
'1' after 25102000 ns, '0' after 25102050 ns,
'1' after 25113000 ns, '0' after 25113050 ns,
'1' after 25124000 ns, '0' after 25124050 ns,
'1' after 25135000 ns, '0' after 25135050 ns,
'1' after 25146000 ns, '0' after 25146050 ns,
'1' after 25157000 ns, '0' after 25157050 ns,
'1' after 25168000 ns, '0' after 25168050 ns,
'1' after 25179000 ns, '0' after 25179050 ns,
'1' after 25190000 ns, '0' after 25190050 ns,
'1' after 25201000 ns, '0' after 25201050 ns,
'1' after 25212000 ns, '0' after 25212050 ns,
'1' after 25223000 ns, '0' after 25223050 ns,
'1' after 25234000 ns, '0' after 25234050 ns,
'1' after 25245000 ns, '0' after 25245050 ns,
'1' after 25256000 ns, '0' after 25256050 ns,
'1' after 25267000 ns, '0' after 25267050 ns,
'1' after 25278000 ns, '0' after 25278050 ns,
'1' after 25289000 ns, '0' after 25289050 ns,
'1' after 25300000 ns, '0' after 25300050 ns,
'1' after 25311000 ns, '0' after 25311050 ns,
'1' after 25322000 ns, '0' after 25322050 ns,
'1' after 25333000 ns, '0' after 25333050 ns,
'1' after 25344000 ns, '0' after 25344050 ns,
'1' after 25355000 ns, '0' after 25355050 ns,
'1' after 25366000 ns, '0' after 25366050 ns,
'1' after 25377000 ns, '0' after 25377050 ns,
'1' after 25388000 ns, '0' after 25388050 ns,
'1' after 25399000 ns, '0' after 25399050 ns,
'1' after 25410000 ns, '0' after 25410050 ns,
'1' after 25421000 ns, '0' after 25421050 ns,
'1' after 25432000 ns, '0' after 25432050 ns,
'1' after 25443000 ns, '0' after 25443050 ns,
'1' after 25454000 ns, '0' after 25454050 ns,
'1' after 25465000 ns, '0' after 25465050 ns,
'1' after 25476000 ns, '0' after 25476050 ns,
'1' after 25487000 ns, '0' after 25487050 ns,
'1' after 25498000 ns, '0' after 25498050 ns,
'1' after 25509000 ns, '0' after 25509050 ns,
'1' after 25520000 ns, '0' after 25520050 ns,
'1' after 25531000 ns, '0' after 25531050 ns,
'1' after 25542000 ns, '0' after 25542050 ns,
'1' after 25553000 ns, '0' after 25553050 ns,
'1' after 25564000 ns, '0' after 25564050 ns,
'1' after 25575000 ns, '0' after 25575050 ns,
'1' after 25586000 ns, '0' after 25586050 ns,
'1' after 25597000 ns, '0' after 25597050 ns,
'1' after 25608000 ns, '0' after 25608050 ns,
'1' after 25619000 ns, '0' after 25619050 ns,
'1' after 25630000 ns, '0' after 25630050 ns,
'1' after 25641000 ns, '0' after 25641050 ns,
'1' after 25652000 ns, '0' after 25652050 ns,
'1' after 25663000 ns, '0' after 25663050 ns,
'1' after 25674000 ns, '0' after 25674050 ns,
'1' after 25685000 ns, '0' after 25685050 ns,
'1' after 25696000 ns, '0' after 25696050 ns,
'1' after 25707000 ns, '0' after 25707050 ns,
'1' after 25718000 ns, '0' after 25718050 ns,
'1' after 25729000 ns, '0' after 25729050 ns,
'1' after 25740000 ns, '0' after 25740050 ns,
'1' after 25751000 ns, '0' after 25751050 ns,
'1' after 25762000 ns, '0' after 25762050 ns,
'1' after 25773000 ns, '0' after 25773050 ns,
'1' after 25784000 ns, '0' after 25784050 ns,
'1' after 25795000 ns, '0' after 25795050 ns,
'1' after 25806000 ns, '0' after 25806050 ns,
'1' after 25817000 ns, '0' after 25817050 ns,
'1' after 25828000 ns, '0' after 25828050 ns,
'1' after 25839000 ns, '0' after 25839050 ns,
'1' after 25850000 ns, '0' after 25850050 ns,
'1' after 25861000 ns, '0' after 25861050 ns,
'1' after 25872000 ns, '0' after 25872050 ns,
'1' after 25883000 ns, '0' after 25883050 ns,
'1' after 25894000 ns, '0' after 25894050 ns,
'1' after 25905000 ns, '0' after 25905050 ns,
'1' after 25916000 ns, '0' after 25916050 ns,
'1' after 25927000 ns, '0' after 25927050 ns,
'1' after 25938000 ns, '0' after 25938050 ns,
'1' after 25949000 ns, '0' after 25949050 ns,
'1' after 25960000 ns, '0' after 25960050 ns,
'1' after 25971000 ns, '0' after 25971050 ns,
'1' after 25982000 ns, '0' after 25982050 ns,
'1' after 25993000 ns, '0' after 25993050 ns,
'1' after 26004000 ns, '0' after 26004050 ns,
'1' after 26015000 ns, '0' after 26015050 ns,
'1' after 26026000 ns, '0' after 26026050 ns,
'1' after 26037000 ns, '0' after 26037050 ns,
'1' after 26048000 ns, '0' after 26048050 ns,
'1' after 26059000 ns, '0' after 26059050 ns,
'1' after 26070000 ns, '0' after 26070050 ns,
'1' after 26081000 ns, '0' after 26081050 ns,
'1' after 26092000 ns, '0' after 26092050 ns,
'1' after 26103000 ns, '0' after 26103050 ns,
'1' after 26114000 ns, '0' after 26114050 ns,
'1' after 26125000 ns, '0' after 26125050 ns,
'1' after 26136000 ns, '0' after 26136050 ns,
'1' after 26147000 ns, '0' after 26147050 ns,
'1' after 26158000 ns, '0' after 26158050 ns,
'1' after 26169000 ns, '0' after 26169050 ns,
'1' after 26180000 ns, '0' after 26180050 ns,
'1' after 26191000 ns, '0' after 26191050 ns,
'1' after 26202000 ns, '0' after 26202050 ns,
'1' after 26213000 ns, '0' after 26213050 ns,
'1' after 26224000 ns, '0' after 26224050 ns,
'1' after 26235000 ns, '0' after 26235050 ns,
'1' after 26246000 ns, '0' after 26246050 ns,
'1' after 26257000 ns, '0' after 26257050 ns,
'1' after 26268000 ns, '0' after 26268050 ns,
'1' after 26279000 ns, '0' after 26279050 ns,
'1' after 26290000 ns, '0' after 26290050 ns,
'1' after 26301000 ns, '0' after 26301050 ns,
'1' after 26312000 ns, '0' after 26312050 ns,
'1' after 26323000 ns, '0' after 26323050 ns,
'1' after 26334000 ns, '0' after 26334050 ns,
'1' after 26345000 ns, '0' after 26345050 ns,
'1' after 26356000 ns, '0' after 26356050 ns,
'1' after 26367000 ns, '0' after 26367050 ns,
'1' after 26378000 ns, '0' after 26378050 ns,
'1' after 26389000 ns, '0' after 26389050 ns,
'1' after 26400000 ns, '0' after 26400050 ns,
'1' after 26411000 ns, '0' after 26411050 ns,
'1' after 26422000 ns, '0' after 26422050 ns,
'1' after 26433000 ns, '0' after 26433050 ns,
'1' after 26444000 ns, '0' after 26444050 ns,
'1' after 26455000 ns, '0' after 26455050 ns,
'1' after 26466000 ns, '0' after 26466050 ns,
'1' after 26477000 ns, '0' after 26477050 ns,
'1' after 26488000 ns, '0' after 26488050 ns,
'1' after 26499000 ns, '0' after 26499050 ns,
'1' after 26510000 ns, '0' after 26510050 ns,
'1' after 26521000 ns, '0' after 26521050 ns,
'1' after 26532000 ns, '0' after 26532050 ns,
'1' after 26543000 ns, '0' after 26543050 ns,
'1' after 26554000 ns, '0' after 26554050 ns,
'1' after 26565000 ns, '0' after 26565050 ns,
'1' after 26576000 ns, '0' after 26576050 ns,
'1' after 26587000 ns, '0' after 26587050 ns,
'1' after 26598000 ns, '0' after 26598050 ns,
'1' after 26609000 ns, '0' after 26609050 ns,
'1' after 26620000 ns, '0' after 26620050 ns,
'1' after 26631000 ns, '0' after 26631050 ns,
'1' after 26642000 ns, '0' after 26642050 ns,
'1' after 26653000 ns, '0' after 26653050 ns,
'1' after 26664000 ns, '0' after 26664050 ns,
'1' after 26675000 ns, '0' after 26675050 ns,
'1' after 26686000 ns, '0' after 26686050 ns,
'1' after 26697000 ns, '0' after 26697050 ns,
'1' after 26708000 ns, '0' after 26708050 ns,
'1' after 26719000 ns, '0' after 26719050 ns,
'1' after 26730000 ns, '0' after 26730050 ns,
'1' after 26741000 ns, '0' after 26741050 ns,
'1' after 26752000 ns, '0' after 26752050 ns,
'1' after 26763000 ns, '0' after 26763050 ns,
'1' after 26774000 ns, '0' after 26774050 ns,
'1' after 26785000 ns, '0' after 26785050 ns,
'1' after 26796000 ns, '0' after 26796050 ns,
'1' after 26807000 ns, '0' after 26807050 ns,
'1' after 26818000 ns, '0' after 26818050 ns,
'1' after 26829000 ns, '0' after 26829050 ns,
'1' after 26840000 ns, '0' after 26840050 ns,
'1' after 26851000 ns, '0' after 26851050 ns,
'1' after 26862000 ns, '0' after 26862050 ns,
'1' after 26873000 ns, '0' after 26873050 ns,
'1' after 26884000 ns, '0' after 26884050 ns,
'1' after 26895000 ns, '0' after 26895050 ns,
'1' after 26906000 ns, '0' after 26906050 ns,
'1' after 26917000 ns, '0' after 26917050 ns,
'1' after 26928000 ns, '0' after 26928050 ns,
'1' after 26939000 ns, '0' after 26939050 ns,
'1' after 26950000 ns, '0' after 26950050 ns,
'1' after 26961000 ns, '0' after 26961050 ns,
'1' after 26972000 ns, '0' after 26972050 ns,
'1' after 26983000 ns, '0' after 26983050 ns,
'1' after 26994000 ns, '0' after 26994050 ns,
'1' after 27005000 ns, '0' after 27005050 ns,
'1' after 27016000 ns, '0' after 27016050 ns,
'1' after 27027000 ns, '0' after 27027050 ns,
'1' after 27038000 ns, '0' after 27038050 ns,
'1' after 27049000 ns, '0' after 27049050 ns,
'1' after 27060000 ns, '0' after 27060050 ns,
'1' after 27071000 ns, '0' after 27071050 ns,
'1' after 27082000 ns, '0' after 27082050 ns,
'1' after 27093000 ns, '0' after 27093050 ns,
'1' after 27104000 ns, '0' after 27104050 ns,
'1' after 27115000 ns, '0' after 27115050 ns,
'1' after 27126000 ns, '0' after 27126050 ns,
'1' after 27137000 ns, '0' after 27137050 ns,
'1' after 27148000 ns, '0' after 27148050 ns,
'1' after 27159000 ns, '0' after 27159050 ns,
'1' after 27170000 ns, '0' after 27170050 ns,
'1' after 27181000 ns, '0' after 27181050 ns,
'1' after 27192000 ns, '0' after 27192050 ns,
'1' after 27203000 ns, '0' after 27203050 ns,
'1' after 27214000 ns, '0' after 27214050 ns,
'1' after 27225000 ns, '0' after 27225050 ns,
'1' after 27236000 ns, '0' after 27236050 ns,
'1' after 27247000 ns, '0' after 27247050 ns,
'1' after 27258000 ns, '0' after 27258050 ns,
'1' after 27269000 ns, '0' after 27269050 ns,
'1' after 27280000 ns, '0' after 27280050 ns,
'1' after 27291000 ns, '0' after 27291050 ns,
'1' after 27302000 ns, '0' after 27302050 ns,
'1' after 27313000 ns, '0' after 27313050 ns,
'1' after 27324000 ns, '0' after 27324050 ns,
'1' after 27335000 ns, '0' after 27335050 ns,
'1' after 27346000 ns, '0' after 27346050 ns,
'1' after 27357000 ns, '0' after 27357050 ns,
'1' after 27368000 ns, '0' after 27368050 ns,
'1' after 27379000 ns, '0' after 27379050 ns,
'1' after 27390000 ns, '0' after 27390050 ns,
'1' after 27401000 ns, '0' after 27401050 ns,
'1' after 27412000 ns, '0' after 27412050 ns,
'1' after 27423000 ns, '0' after 27423050 ns,
'1' after 27434000 ns, '0' after 27434050 ns,
'1' after 27445000 ns, '0' after 27445050 ns,
'1' after 27456000 ns, '0' after 27456050 ns,
'1' after 27467000 ns, '0' after 27467050 ns,
'1' after 27478000 ns, '0' after 27478050 ns,
'1' after 27489000 ns, '0' after 27489050 ns,
'1' after 27500000 ns, '0' after 27500050 ns,
'1' after 27511000 ns, '0' after 27511050 ns,
'1' after 27522000 ns, '0' after 27522050 ns,
'1' after 27533000 ns, '0' after 27533050 ns,
'1' after 27544000 ns, '0' after 27544050 ns,
'1' after 27555000 ns, '0' after 27555050 ns,
'1' after 27566000 ns, '0' after 27566050 ns,
'1' after 27577000 ns, '0' after 27577050 ns,
'1' after 27588000 ns, '0' after 27588050 ns,
'1' after 27599000 ns, '0' after 27599050 ns,
'1' after 27610000 ns, '0' after 27610050 ns,
'1' after 27621000 ns, '0' after 27621050 ns,
'1' after 27632000 ns, '0' after 27632050 ns,
'1' after 27643000 ns, '0' after 27643050 ns,
'1' after 27654000 ns, '0' after 27654050 ns,
'1' after 27665000 ns, '0' after 27665050 ns,
'1' after 27676000 ns, '0' after 27676050 ns,
'1' after 27687000 ns, '0' after 27687050 ns,
'1' after 27698000 ns, '0' after 27698050 ns,
'1' after 27709000 ns, '0' after 27709050 ns,
'1' after 27720000 ns, '0' after 27720050 ns,
'1' after 27731000 ns, '0' after 27731050 ns,
'1' after 27742000 ns, '0' after 27742050 ns,
'1' after 27753000 ns, '0' after 27753050 ns,
'1' after 27764000 ns, '0' after 27764050 ns,
'1' after 27775000 ns, '0' after 27775050 ns,
'1' after 27786000 ns, '0' after 27786050 ns,
'1' after 27797000 ns, '0' after 27797050 ns,
'1' after 27808000 ns, '0' after 27808050 ns,
'1' after 27819000 ns, '0' after 27819050 ns,
'1' after 27830000 ns, '0' after 27830050 ns,
'1' after 27841000 ns, '0' after 27841050 ns,
'1' after 27852000 ns, '0' after 27852050 ns,
'1' after 27863000 ns, '0' after 27863050 ns,
'1' after 27874000 ns, '0' after 27874050 ns,
'1' after 27885000 ns, '0' after 27885050 ns,
'1' after 27896000 ns, '0' after 27896050 ns,
'1' after 27907000 ns, '0' after 27907050 ns,
'1' after 27918000 ns, '0' after 27918050 ns,
'1' after 27929000 ns, '0' after 27929050 ns,
'1' after 27940000 ns, '0' after 27940050 ns,
'1' after 27951000 ns, '0' after 27951050 ns,
'1' after 27962000 ns, '0' after 27962050 ns,
'1' after 27973000 ns, '0' after 27973050 ns,
'1' after 27984000 ns, '0' after 27984050 ns,
'1' after 27995000 ns, '0' after 27995050 ns,
'1' after 28006000 ns, '0' after 28006050 ns,
'1' after 28017000 ns, '0' after 28017050 ns,
'1' after 28028000 ns, '0' after 28028050 ns,
'1' after 28039000 ns, '0' after 28039050 ns,
'1' after 28050000 ns, '0' after 28050050 ns,
'1' after 28061000 ns, '0' after 28061050 ns,
'1' after 28072000 ns, '0' after 28072050 ns,
'1' after 28083000 ns, '0' after 28083050 ns,
'1' after 28094000 ns, '0' after 28094050 ns,
'1' after 28105000 ns, '0' after 28105050 ns,
'1' after 28116000 ns, '0' after 28116050 ns,
'1' after 28127000 ns, '0' after 28127050 ns,
'1' after 28138000 ns, '0' after 28138050 ns,
'1' after 28149000 ns, '0' after 28149050 ns,
'1' after 28160000 ns, '0' after 28160050 ns,
'1' after 28171000 ns, '0' after 28171050 ns,
'1' after 28182000 ns, '0' after 28182050 ns,
'1' after 28193000 ns, '0' after 28193050 ns,
'1' after 28204000 ns, '0' after 28204050 ns,
'1' after 28215000 ns, '0' after 28215050 ns,
'1' after 28226000 ns, '0' after 28226050 ns,
'1' after 28237000 ns, '0' after 28237050 ns,
'1' after 28248000 ns, '0' after 28248050 ns,
'1' after 28259000 ns, '0' after 28259050 ns,
'1' after 28270000 ns, '0' after 28270050 ns,
'1' after 28281000 ns, '0' after 28281050 ns,
'1' after 28292000 ns, '0' after 28292050 ns,
'1' after 28303000 ns, '0' after 28303050 ns,
'1' after 28314000 ns, '0' after 28314050 ns,
'1' after 28325000 ns, '0' after 28325050 ns,
'1' after 28336000 ns, '0' after 28336050 ns,
'1' after 28347000 ns, '0' after 28347050 ns,
'1' after 28358000 ns, '0' after 28358050 ns,
'1' after 28369000 ns, '0' after 28369050 ns,
'1' after 28380000 ns, '0' after 28380050 ns,
'1' after 28391000 ns, '0' after 28391050 ns,
'1' after 28402000 ns, '0' after 28402050 ns,
'1' after 28413000 ns, '0' after 28413050 ns,
'1' after 28424000 ns, '0' after 28424050 ns,
'1' after 28435000 ns, '0' after 28435050 ns,
'1' after 28446000 ns, '0' after 28446050 ns,
'1' after 28457000 ns, '0' after 28457050 ns,
'1' after 28468000 ns, '0' after 28468050 ns,
'1' after 28479000 ns, '0' after 28479050 ns,
'1' after 28490000 ns, '0' after 28490050 ns,
'1' after 28501000 ns, '0' after 28501050 ns,
'1' after 28512000 ns, '0' after 28512050 ns,
'1' after 28523000 ns, '0' after 28523050 ns,
'1' after 28534000 ns, '0' after 28534050 ns,
'1' after 28545000 ns, '0' after 28545050 ns,
'1' after 28556000 ns, '0' after 28556050 ns,
'1' after 28567000 ns, '0' after 28567050 ns,
'1' after 28578000 ns, '0' after 28578050 ns,
'1' after 28589000 ns, '0' after 28589050 ns,
'1' after 28600000 ns, '0' after 28600050 ns,
'1' after 28611000 ns, '0' after 28611050 ns,
'1' after 28622000 ns, '0' after 28622050 ns,
'1' after 28633000 ns, '0' after 28633050 ns,
'1' after 28644000 ns, '0' after 28644050 ns,
'1' after 28655000 ns, '0' after 28655050 ns,
'1' after 28666000 ns, '0' after 28666050 ns,
'1' after 28677000 ns, '0' after 28677050 ns,
'1' after 28688000 ns, '0' after 28688050 ns,
'1' after 28699000 ns, '0' after 28699050 ns,
'1' after 28710000 ns, '0' after 28710050 ns,
'1' after 28721000 ns, '0' after 28721050 ns,
'1' after 28732000 ns, '0' after 28732050 ns,
'1' after 28743000 ns, '0' after 28743050 ns,
'1' after 28754000 ns, '0' after 28754050 ns,
'1' after 28765000 ns, '0' after 28765050 ns,
'1' after 28776000 ns, '0' after 28776050 ns,
'1' after 28787000 ns, '0' after 28787050 ns,
'1' after 28798000 ns, '0' after 28798050 ns,
'1' after 28809000 ns, '0' after 28809050 ns,
'1' after 28820000 ns, '0' after 28820050 ns,
'1' after 28831000 ns, '0' after 28831050 ns,
'1' after 28842000 ns, '0' after 28842050 ns,
'1' after 28853000 ns, '0' after 28853050 ns,
'1' after 28864000 ns, '0' after 28864050 ns,
'1' after 28875000 ns, '0' after 28875050 ns,
'1' after 28886000 ns, '0' after 28886050 ns,
'1' after 28897000 ns, '0' after 28897050 ns,
'1' after 28908000 ns, '0' after 28908050 ns,
'1' after 28919000 ns, '0' after 28919050 ns,
'1' after 28930000 ns, '0' after 28930050 ns,
'1' after 28941000 ns, '0' after 28941050 ns,
'1' after 28952000 ns, '0' after 28952050 ns,
'1' after 28963000 ns, '0' after 28963050 ns,
'1' after 28974000 ns, '0' after 28974050 ns,
'1' after 28985000 ns, '0' after 28985050 ns,
'1' after 28996000 ns, '0' after 28996050 ns,
'1' after 29007000 ns, '0' after 29007050 ns,
'1' after 29018000 ns, '0' after 29018050 ns,
'1' after 29029000 ns, '0' after 29029050 ns,
'1' after 29040000 ns, '0' after 29040050 ns,
'1' after 29051000 ns, '0' after 29051050 ns,
'1' after 29062000 ns, '0' after 29062050 ns,
'1' after 29073000 ns, '0' after 29073050 ns,
'1' after 29084000 ns, '0' after 29084050 ns,
'1' after 29095000 ns, '0' after 29095050 ns,
'1' after 29106000 ns, '0' after 29106050 ns,
'1' after 29117000 ns, '0' after 29117050 ns,
'1' after 29128000 ns, '0' after 29128050 ns,
'1' after 29139000 ns, '0' after 29139050 ns,
'1' after 29150000 ns, '0' after 29150050 ns,
'1' after 29161000 ns, '0' after 29161050 ns,
'1' after 29172000 ns, '0' after 29172050 ns,
'1' after 29183000 ns, '0' after 29183050 ns,
'1' after 29194000 ns, '0' after 29194050 ns,
'1' after 29205000 ns, '0' after 29205050 ns,
'1' after 29216000 ns, '0' after 29216050 ns,
'1' after 29227000 ns, '0' after 29227050 ns,
'1' after 29238000 ns, '0' after 29238050 ns,
'1' after 29249000 ns, '0' after 29249050 ns,
'1' after 29260000 ns, '0' after 29260050 ns,
'1' after 29271000 ns, '0' after 29271050 ns,
'1' after 29282000 ns, '0' after 29282050 ns,
'1' after 29293000 ns, '0' after 29293050 ns,
'1' after 29304000 ns, '0' after 29304050 ns,
'1' after 29315000 ns, '0' after 29315050 ns,
'1' after 29326000 ns, '0' after 29326050 ns,
'1' after 29337000 ns, '0' after 29337050 ns,
'1' after 29348000 ns, '0' after 29348050 ns;

 -- intr_sig <= '0', '1' after 1000 ns, '0' after 1050 ns;
 -- port_io_sig(30 downto 27) <= "0000", "1000" after 8000 ns;
  --port_io_sig(3 downto 0) <= "1111";
  port_io_sig(29 downto 0) <= (others => 'Z');
  port_io_sig(31) <= '0', '1' after 31803511 ns, '0' after 31803611 ns;
  port_io_sig(30) <= '0';

end architecture behavior;
