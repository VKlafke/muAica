library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.muAica_pkg.all;

entity muAica_tb is
end entity muAica_tb;

architecture behavior of muAica_tb is

  -- processor top module component
  COMPONENT muAica is
    port (
      clk       : in    std_logic;
      rst_bt    : in    std_logic;
      port_io   : inout std_logic_vector (n-1 downto 0); -- configurable IO port
      tx        : out std_logic;
	    rx: in std_logic
    );
  end COMPONENT muAica;

  -- System clock and reset
  signal  clk   : std_logic;
  signal  rst_bt: std_logic;

  constant half_period : time := 10 ns; -- 50 MHZ

  signal  intr_sig : std_logic;
  signal  port_io_sig  : std_logic_vector (n-1 downto 0); -- interface with microcontroller port

  signal tx_s : std_logic; -- tx signal
  signal rx_s : std_logic;

  signal tx_dv : std_logic;
  signal tx_active_s : std_logic;
  signal tx_done :std_logic;
  signal data_tx : std_logic_vector(7 downto 0);

begin

  -- Clock process: 100 MHz
  signal_clk : process
  begin
    clk <= '0'; wait for half_period;
    loop
      clk <= '1'; wait for half_period;
      clk <= '0'; wait for half_period;
    end loop;
  end process signal_clk;

  -- Clock
  rst_button : process -- debounce should be disabled inside 'aica/bt_debounce' (stability time ~0)
  begin
    rst_bt <= '0'; wait for 100 ns;
    loop
      rst_bt <= '1'; wait for 50 ns;
      rst_bt <= '0'; wait for 20 sec;
      rst_bt <= '1'; wait for 100 ns;
      rst_bt <= '0'; wait for 10 sec;
    end loop;
  end process rst_button;

-- Port Map
  MICRO_AICA: muAica
  port map(
    clk     => clk,
    rst_bt  => rst_bt,
    port_io => port_io_sig,
    tx      => tx_s,
	  rx		=> rx_s
  );
  
 -- rx_s <= '0';

  -- Send data to rx
  TX_DATA_SEND: entity work.UART_TX_v1
  port map(
    i_Clk       => clk,
    i_TX_DV     => tx_dv,
    i_TX_Byte   => data_tx,
    o_TX_Active => tx_active_s,
    o_TX_Serial => rx_s,
    o_TX_Done   => tx_done
  );

  -- VHDL for data_tx:
data_tx <= x"00" after 0 ns,
x"00" after 10850 ns,
x"07" after 21700 ns,
x"70" after 32550 ns,
x"17" after 43400 ns,
x"21" after 54250 ns,
x"00" after 65100 ns,
x"00" after 75950 ns,
x"13" after 86800 ns,
x"01" after 97650 ns,
x"41" after 108500 ns,
x"56" after 119350 ns,
x"13" after 130200 ns,
x"01" after 141050 ns,
x"C1" after 151900 ns,
x"FF" after 162750 ns,
x"23" after 173600 ns,
x"20" after 184450 ns,
x"11" after 195300 ns,
x"00" after 206150 ns,
x"37" after 217000 ns,
x"1F" after 227850 ns,
x"00" after 238700 ns,
x"00" after 249550 ns,
x"13" after 260400 ns,
x"0F" after 271250 ns,
x"0F" after 282100 ns,
x"80" after 292950 ns,
x"73" after 303800 ns,
x"20" after 314650 ns,
x"4F" after 325500 ns,
x"30" after 336350 ns,
x"73" after 347200 ns,
x"60" after 358050 ns,
x"44" after 368900 ns,
x"30" after 379750 ns,
x"73" after 390600 ns,
x"60" after 401450 ns,
x"04" after 412300 ns,
x"30" after 423150 ns,
x"73" after 434000 ns,
x"10" after 444850 ns,
x"10" after 455700 ns,
x"34" after 466550 ns,
x"73" after 477400 ns,
x"10" after 488250 ns,
x"20" after 499100 ns,
x"34" after 509950 ns,
x"EF" after 520800 ns,
x"00" after 531650 ns,
x"00" after 542500 ns,
x"6C" after 553350 ns,
x"83" after 564200 ns,
x"20" after 575050 ns,
x"01" after 585900 ns,
x"00" after 596750 ns,
x"13" after 607600 ns,
x"01" after 618450 ns,
x"41" after 629300 ns,
x"00" after 640150 ns,
x"67" after 651000 ns,
x"80" after 661850 ns,
x"00" after 672700 ns,
x"00" after 683550 ns,
x"93" after 694400 ns,
x"08" after 705250 ns,
x"10" after 716100 ns,
x"00" after 726950 ns,
x"73" after 737800 ns,
x"00" after 748650 ns,
x"00" after 759500 ns,
x"00" after 770350 ns,
x"67" after 781200 ns,
x"80" after 792050 ns,
x"00" after 802900 ns,
x"00" after 813750 ns,
x"93" after 824600 ns,
x"08" after 835450 ns,
x"20" after 846300 ns,
x"00" after 857150 ns,
x"73" after 868000 ns,
x"00" after 878850 ns,
x"00" after 889700 ns,
x"00" after 900550 ns,
x"67" after 911400 ns,
x"80" after 922250 ns,
x"00" after 933100 ns,
x"00" after 943950 ns,
x"93" after 954800 ns,
x"08" after 965650 ns,
x"30" after 976500 ns,
x"00" after 987350 ns,
x"73" after 998200 ns,
x"00" after 1009050 ns,
x"00" after 1019900 ns,
x"00" after 1030750 ns,
x"67" after 1041600 ns,
x"80" after 1052450 ns,
x"00" after 1063300 ns,
x"00" after 1074150 ns,
x"93" after 1085000 ns,
x"08" after 1095850 ns,
x"40" after 1106700 ns,
x"00" after 1117550 ns,
x"73" after 1128400 ns,
x"00" after 1139250 ns,
x"00" after 1150100 ns,
x"00" after 1160950 ns,
x"67" after 1171800 ns,
x"80" after 1182650 ns,
x"00" after 1193500 ns,
x"00" after 1204350 ns,
x"93" after 1215200 ns,
x"08" after 1226050 ns,
x"A0" after 1236900 ns,
x"00" after 1247750 ns,
x"73" after 1258600 ns,
x"00" after 1269450 ns,
x"00" after 1280300 ns,
x"00" after 1291150 ns,
x"67" after 1302000 ns,
x"80" after 1312850 ns,
x"00" after 1323700 ns,
x"00" after 1334550 ns,
x"93" after 1345400 ns,
x"08" after 1356250 ns,
x"B0" after 1367100 ns,
x"00" after 1377950 ns,
x"73" after 1388800 ns,
x"00" after 1399650 ns,
x"00" after 1410500 ns,
x"00" after 1421350 ns,
x"67" after 1432200 ns,
x"80" after 1443050 ns,
x"00" after 1453900 ns,
x"00" after 1464750 ns,
x"93" after 1475600 ns,
x"08" after 1486450 ns,
x"C0" after 1497300 ns,
x"00" after 1508150 ns,
x"73" after 1519000 ns,
x"00" after 1529850 ns,
x"00" after 1540700 ns,
x"00" after 1551550 ns,
x"67" after 1562400 ns,
x"80" after 1573250 ns,
x"00" after 1584100 ns,
x"00" after 1594950 ns,
x"93" after 1605800 ns,
x"08" after 1616650 ns,
x"D0" after 1627500 ns,
x"00" after 1638350 ns,
x"73" after 1649200 ns,
x"00" after 1660050 ns,
x"00" after 1670900 ns,
x"00" after 1681750 ns,
x"67" after 1692600 ns,
x"80" after 1703450 ns,
x"00" after 1714300 ns,
x"00" after 1725150 ns,
x"93" after 1736000 ns,
x"08" after 1746850 ns,
x"E0" after 1757700 ns,
x"00" after 1768550 ns,
x"73" after 1779400 ns,
x"00" after 1790250 ns,
x"00" after 1801100 ns,
x"00" after 1811950 ns,
x"67" after 1822800 ns,
x"80" after 1833650 ns,
x"00" after 1844500 ns,
x"00" after 1855350 ns,
x"93" after 1866200 ns,
x"08" after 1877050 ns,
x"F0" after 1887900 ns,
x"00" after 1898750 ns,
x"73" after 1909600 ns,
x"00" after 1920450 ns,
x"00" after 1931300 ns,
x"00" after 1942150 ns,
x"67" after 1953000 ns,
x"80" after 1963850 ns,
x"00" after 1974700 ns,
x"00" after 1985550 ns,
x"13" after 1996400 ns,
x"01" after 2007250 ns,
x"81" after 2018100 ns,
x"FE" after 2028950 ns,
x"23" after 2039800 ns,
x"2A" after 2050650 ns,
x"81" after 2061500 ns,
x"00" after 2072350 ns,
x"13" after 2083200 ns,
x"04" after 2094050 ns,
x"81" after 2104900 ns,
x"01" after 2115750 ns,
x"23" after 2126600 ns,
x"26" after 2137450 ns,
x"A4" after 2148300 ns,
x"FE" after 2159150 ns,
x"83" after 2170000 ns,
x"27" after 2180850 ns,
x"C4" after 2191700 ns,
x"FE" after 2202550 ns,
x"23" after 2213400 ns,
x"2A" after 2224250 ns,
x"F4" after 2235100 ns,
x"FE" after 2245950 ns,
x"6F" after 2256800 ns,
x"00" after 2267650 ns,
x"00" after 2278500 ns,
x"01" after 2289350 ns,
x"83" after 2300200 ns,
x"27" after 2311050 ns,
x"44" after 2321900 ns,
x"FF" after 2332750 ns,
x"93" after 2343600 ns,
x"87" after 2354450 ns,
x"17" after 2365300 ns,
x"00" after 2376150 ns,
x"23" after 2387000 ns,
x"2A" after 2397850 ns,
x"F4" after 2408700 ns,
x"FE" after 2419550 ns,
x"83" after 2430400 ns,
x"27" after 2441250 ns,
x"44" after 2452100 ns,
x"FF" after 2462950 ns,
x"83" after 2473800 ns,
x"C7" after 2484650 ns,
x"07" after 2495500 ns,
x"00" after 2506350 ns,
x"E3" after 2517200 ns,
x"96" after 2528050 ns,
x"07" after 2538900 ns,
x"FE" after 2549750 ns,
x"03" after 2560600 ns,
x"27" after 2571450 ns,
x"44" after 2582300 ns,
x"FF" after 2593150 ns,
x"83" after 2604000 ns,
x"27" after 2614850 ns,
x"C4" after 2625700 ns,
x"FE" after 2636550 ns,
x"B3" after 2647400 ns,
x"07" after 2658250 ns,
x"F7" after 2669100 ns,
x"40" after 2679950 ns,
x"13" after 2690800 ns,
x"85" after 2701650 ns,
x"07" after 2712500 ns,
x"00" after 2723350 ns,
x"03" after 2734200 ns,
x"24" after 2745050 ns,
x"41" after 2755900 ns,
x"01" after 2766750 ns,
x"13" after 2777600 ns,
x"01" after 2788450 ns,
x"81" after 2799300 ns,
x"01" after 2810150 ns,
x"67" after 2821000 ns,
x"80" after 2831850 ns,
x"00" after 2842700 ns,
x"00" after 2853550 ns,
x"13" after 2864400 ns,
x"01" after 2875250 ns,
x"81" after 2886100 ns,
x"FE" after 2896950 ns,
x"23" after 2907800 ns,
x"2A" after 2918650 ns,
x"81" after 2929500 ns,
x"00" after 2940350 ns,
x"13" after 2951200 ns,
x"04" after 2962050 ns,
x"81" after 2972900 ns,
x"01" after 2983750 ns,
x"23" after 2994600 ns,
x"26" after 3005450 ns,
x"A4" after 3016300 ns,
x"FE" after 3027150 ns,
x"23" after 3038000 ns,
x"24" after 3048850 ns,
x"B4" after 3059700 ns,
x"FE" after 3070550 ns,
x"23" after 3081400 ns,
x"2A" after 3092250 ns,
x"04" after 3103100 ns,
x"FE" after 3113950 ns,
x"6F" after 3124800 ns,
x"00" after 3135650 ns,
x"00" after 3146500 ns,
x"03" after 3157350 ns,
x"03" after 3168200 ns,
x"27" after 3179050 ns,
x"84" after 3189900 ns,
x"FE" after 3200750 ns,
x"93" after 3211600 ns,
x"07" after 3222450 ns,
x"17" after 3233300 ns,
x"00" after 3244150 ns,
x"23" after 3255000 ns,
x"24" after 3265850 ns,
x"F4" after 3276700 ns,
x"FE" after 3287550 ns,
x"83" after 3298400 ns,
x"27" after 3309250 ns,
x"C4" after 3320100 ns,
x"FE" after 3330950 ns,
x"93" after 3341800 ns,
x"86" after 3352650 ns,
x"17" after 3363500 ns,
x"00" after 3374350 ns,
x"23" after 3385200 ns,
x"26" after 3396050 ns,
x"D4" after 3406900 ns,
x"FE" after 3417750 ns,
x"03" after 3428600 ns,
x"47" after 3439450 ns,
x"07" after 3450300 ns,
x"00" after 3461150 ns,
x"23" after 3472000 ns,
x"80" after 3482850 ns,
x"E7" after 3493700 ns,
x"00" after 3504550 ns,
x"83" after 3515400 ns,
x"27" after 3526250 ns,
x"44" after 3537100 ns,
x"FF" after 3547950 ns,
x"93" after 3558800 ns,
x"87" after 3569650 ns,
x"17" after 3580500 ns,
x"00" after 3591350 ns,
x"23" after 3602200 ns,
x"2A" after 3613050 ns,
x"F4" after 3623900 ns,
x"FE" after 3634750 ns,
x"83" after 3645600 ns,
x"27" after 3656450 ns,
x"84" after 3667300 ns,
x"FE" after 3678150 ns,
x"83" after 3689000 ns,
x"C7" after 3699850 ns,
x"07" after 3710700 ns,
x"00" after 3721550 ns,
x"E3" after 3732400 ns,
x"96" after 3743250 ns,
x"07" after 3754100 ns,
x"FC" after 3764950 ns,
x"83" after 3775800 ns,
x"27" after 3786650 ns,
x"C4" after 3797500 ns,
x"FE" after 3808350 ns,
x"23" after 3819200 ns,
x"80" after 3830050 ns,
x"07" after 3840900 ns,
x"00" after 3851750 ns,
x"83" after 3862600 ns,
x"27" after 3873450 ns,
x"44" after 3884300 ns,
x"FF" after 3895150 ns,
x"13" after 3906000 ns,
x"85" after 3916850 ns,
x"07" after 3927700 ns,
x"00" after 3938550 ns,
x"03" after 3949400 ns,
x"24" after 3960250 ns,
x"41" after 3971100 ns,
x"01" after 3981950 ns,
x"13" after 3992800 ns,
x"01" after 4003650 ns,
x"81" after 4014500 ns,
x"01" after 4025350 ns,
x"67" after 4036200 ns,
x"80" after 4047050 ns,
x"00" after 4057900 ns,
x"00" after 4068750 ns,
x"13" after 4079600 ns,
x"01" after 4090450 ns,
x"81" after 4101300 ns,
x"FD" after 4112150 ns,
x"23" after 4123000 ns,
x"22" after 4133850 ns,
x"81" after 4144700 ns,
x"02" after 4155550 ns,
x"13" after 4166400 ns,
x"04" after 4177250 ns,
x"81" after 4188100 ns,
x"02" after 4198950 ns,
x"23" after 4209800 ns,
x"2E" after 4220650 ns,
x"A4" after 4231500 ns,
x"FC" after 4242350 ns,
x"23" after 4253200 ns,
x"2C" after 4264050 ns,
x"B4" after 4274900 ns,
x"FC" after 4285750 ns,
x"B7" after 4296600 ns,
x"17" after 4307450 ns,
x"00" after 4318300 ns,
x"00" after 4329150 ns,
x"93" after 4340000 ns,
x"87" after 4350850 ns,
x"87" after 4361700 ns,
x"80" after 4372550 ns,
x"83" after 4383400 ns,
x"A5" after 4394250 ns,
x"07" after 4405100 ns,
x"00" after 4415950 ns,
x"03" after 4426800 ns,
x"A6" after 4437650 ns,
x"47" after 4448500 ns,
x"00" after 4459350 ns,
x"83" after 4470200 ns,
x"A6" after 4481050 ns,
x"87" after 4491900 ns,
x"00" after 4502750 ns,
x"03" after 4513600 ns,
x"A7" after 4524450 ns,
x"C7" after 4535300 ns,
x"00" after 4546150 ns,
x"23" after 4557000 ns,
x"22" after 4567850 ns,
x"B4" after 4578700 ns,
x"FE" after 4589550 ns,
x"23" after 4600400 ns,
x"24" after 4611250 ns,
x"C4" after 4622100 ns,
x"FE" after 4632950 ns,
x"23" after 4643800 ns,
x"26" after 4654650 ns,
x"D4" after 4665500 ns,
x"FE" after 4676350 ns,
x"23" after 4687200 ns,
x"28" after 4698050 ns,
x"E4" after 4708900 ns,
x"FE" after 4719750 ns,
x"83" after 4730600 ns,
x"C7" after 4741450 ns,
x"07" after 4752300 ns,
x"01" after 4763150 ns,
x"23" after 4774000 ns,
x"0A" after 4784850 ns,
x"F4" after 4795700 ns,
x"FE" after 4806550 ns,
x"83" after 4817400 ns,
x"27" after 4828250 ns,
x"84" after 4839100 ns,
x"FD" after 4849950 ns,
x"93" after 4860800 ns,
x"D7" after 4871650 ns,
x"47" after 4882500 ns,
x"40" after 4893350 ns,
x"93" after 4904200 ns,
x"F7" after 4915050 ns,
x"F7" after 4925900 ns,
x"00" after 4936750 ns,
x"93" after 4947600 ns,
x"87" after 4958450 ns,
x"87" after 4969300 ns,
x"FF" after 4980150 ns,
x"B3" after 4991000 ns,
x"87" after 5001850 ns,
x"87" after 5012700 ns,
x"00" after 5023550 ns,
x"03" after 5034400 ns,
x"C7" after 5045250 ns,
x"C7" after 5056100 ns,
x"FE" after 5066950 ns,
x"83" after 5077800 ns,
x"27" after 5088650 ns,
x"C4" after 5099500 ns,
x"FD" after 5110350 ns,
x"23" after 5121200 ns,
x"80" after 5132050 ns,
x"E7" after 5142900 ns,
x"00" after 5153750 ns,
x"83" after 5164600 ns,
x"27" after 5175450 ns,
x"84" after 5186300 ns,
x"FD" after 5197150 ns,
x"13" after 5208000 ns,
x"F7" after 5218850 ns,
x"F7" after 5229700 ns,
x"00" after 5240550 ns,
x"83" after 5251400 ns,
x"27" after 5262250 ns,
x"C4" after 5273100 ns,
x"FD" after 5283950 ns,
x"93" after 5294800 ns,
x"87" after 5305650 ns,
x"17" after 5316500 ns,
x"00" after 5327350 ns,
x"13" after 5338200 ns,
x"07" after 5349050 ns,
x"87" after 5359900 ns,
x"FF" after 5370750 ns,
x"33" after 5381600 ns,
x"07" after 5392450 ns,
x"87" after 5403300 ns,
x"00" after 5414150 ns,
x"03" after 5425000 ns,
x"47" after 5435850 ns,
x"C7" after 5446700 ns,
x"FE" after 5457550 ns,
x"23" after 5468400 ns,
x"80" after 5479250 ns,
x"E7" after 5490100 ns,
x"00" after 5500950 ns,
x"83" after 5511800 ns,
x"27" after 5522650 ns,
x"C4" after 5533500 ns,
x"FD" after 5544350 ns,
x"93" after 5555200 ns,
x"87" after 5566050 ns,
x"27" after 5576900 ns,
x"00" after 5587750 ns,
x"23" after 5598600 ns,
x"80" after 5609450 ns,
x"07" after 5620300 ns,
x"00" after 5631150 ns,
x"93" after 5642000 ns,
x"07" after 5652850 ns,
x"20" after 5663700 ns,
x"00" after 5674550 ns,
x"13" after 5685400 ns,
x"85" after 5696250 ns,
x"07" after 5707100 ns,
x"00" after 5717950 ns,
x"03" after 5728800 ns,
x"24" after 5739650 ns,
x"41" after 5750500 ns,
x"02" after 5761350 ns,
x"13" after 5772200 ns,
x"01" after 5783050 ns,
x"81" after 5793900 ns,
x"02" after 5804750 ns,
x"67" after 5815600 ns,
x"80" after 5826450 ns,
x"00" after 5837300 ns,
x"00" after 5848150 ns,
x"13" after 5859000 ns,
x"01" after 5869850 ns,
x"01" after 5880700 ns,
x"FC" after 5891550 ns,
x"23" after 5902400 ns,
x"2E" after 5913250 ns,
x"81" after 5924100 ns,
x"02" after 5934950 ns,
x"13" after 5945800 ns,
x"04" after 5956650 ns,
x"01" after 5967500 ns,
x"04" after 5978350 ns,
x"23" after 5989200 ns,
x"22" after 6000050 ns,
x"A4" after 6010900 ns,
x"FC" after 6021750 ns,
x"23" after 6032600 ns,
x"20" after 6043450 ns,
x"B4" after 6054300 ns,
x"FC" after 6065150 ns,
x"23" after 6076000 ns,
x"2A" after 6086850 ns,
x"04" after 6097700 ns,
x"FE" after 6108550 ns,
x"23" after 6119400 ns,
x"26" after 6130250 ns,
x"04" after 6141100 ns,
x"FE" after 6151950 ns,
x"83" after 6162800 ns,
x"27" after 6173650 ns,
x"04" after 6184500 ns,
x"FC" after 6195350 ns,
x"93" after 6206200 ns,
x"D7" after 6217050 ns,
x"F7" after 6227900 ns,
x"01" after 6238750 ns,
x"93" after 6249600 ns,
x"F7" after 6260450 ns,
x"F7" after 6271300 ns,
x"0F" after 6282150 ns,
x"23" after 6293000 ns,
x"24" after 6303850 ns,
x"F4" after 6314700 ns,
x"FE" after 6325550 ns,
x"83" after 6336400 ns,
x"27" after 6347250 ns,
x"84" after 6358100 ns,
x"FE" after 6368950 ns,
x"63" after 6379800 ns,
x"88" after 6390650 ns,
x"07" after 6401500 ns,
x"00" after 6412350 ns,
x"83" after 6423200 ns,
x"27" after 6434050 ns,
x"04" after 6444900 ns,
x"FC" after 6455750 ns,
x"B3" after 6466600 ns,
x"07" after 6477450 ns,
x"F0" after 6488300 ns,
x"40" after 6499150 ns,
x"23" after 6510000 ns,
x"20" after 6520850 ns,
x"F4" after 6531700 ns,
x"FC" after 6542550 ns,
x"03" after 6553400 ns,
x"27" after 6564250 ns,
x"04" after 6575100 ns,
x"FC" after 6585950 ns,
x"93" after 6596800 ns,
x"07" after 6607650 ns,
x"A0" after 6618500 ns,
x"00" after 6629350 ns,
x"B3" after 6640200 ns,
x"67" after 6651050 ns,
x"F7" after 6661900 ns,
x"02" after 6672750 ns,
x"13" after 6683600 ns,
x"F7" after 6694450 ns,
x"F7" after 6705300 ns,
x"0F" after 6716150 ns,
x"83" after 6727000 ns,
x"27" after 6737850 ns,
x"44" after 6748700 ns,
x"FF" after 6759550 ns,
x"93" after 6770400 ns,
x"86" after 6781250 ns,
x"17" after 6792100 ns,
x"00" after 6802950 ns,
x"23" after 6813800 ns,
x"2A" after 6824650 ns,
x"D4" after 6835500 ns,
x"FE" after 6846350 ns,
x"13" after 6857200 ns,
x"07" after 6868050 ns,
x"07" after 6878900 ns,
x"03" after 6889750 ns,
x"13" after 6900600 ns,
x"77" after 6911450 ns,
x"F7" after 6922300 ns,
x"0F" after 6933150 ns,
x"93" after 6944000 ns,
x"87" after 6954850 ns,
x"87" after 6965700 ns,
x"FF" after 6976550 ns,
x"B3" after 6987400 ns,
x"87" after 6998250 ns,
x"87" after 7009100 ns,
x"00" after 7019950 ns,
x"23" after 7030800 ns,
x"88" after 7041650 ns,
x"E7" after 7052500 ns,
x"FC" after 7063350 ns,
x"03" after 7074200 ns,
x"27" after 7085050 ns,
x"04" after 7095900 ns,
x"FC" after 7106750 ns,
x"93" after 7117600 ns,
x"07" after 7128450 ns,
x"A0" after 7139300 ns,
x"00" after 7150150 ns,
x"B3" after 7161000 ns,
x"47" after 7171850 ns,
x"F7" after 7182700 ns,
x"02" after 7193550 ns,
x"23" after 7204400 ns,
x"20" after 7215250 ns,
x"F4" after 7226100 ns,
x"FC" after 7236950 ns,
x"83" after 7247800 ns,
x"27" after 7258650 ns,
x"04" after 7269500 ns,
x"FC" after 7280350 ns,
x"E3" after 7291200 ns,
x"9E" after 7302050 ns,
x"07" after 7312900 ns,
x"FA" after 7323750 ns,
x"83" after 7334600 ns,
x"27" after 7345450 ns,
x"84" after 7356300 ns,
x"FE" after 7367150 ns,
x"63" after 7378000 ns,
x"80" after 7388850 ns,
x"07" after 7399700 ns,
x"02" after 7410550 ns,
x"83" after 7421400 ns,
x"27" after 7432250 ns,
x"44" after 7443100 ns,
x"FF" after 7453950 ns,
x"13" after 7464800 ns,
x"87" after 7475650 ns,
x"17" after 7486500 ns,
x"00" after 7497350 ns,
x"23" after 7508200 ns,
x"2A" after 7519050 ns,
x"E4" after 7529900 ns,
x"FE" after 7540750 ns,
x"93" after 7551600 ns,
x"87" after 7562450 ns,
x"87" after 7573300 ns,
x"FF" after 7584150 ns,
x"B3" after 7595000 ns,
x"87" after 7605850 ns,
x"87" after 7616700 ns,
x"00" after 7627550 ns,
x"13" after 7638400 ns,
x"07" after 7649250 ns,
x"D0" after 7660100 ns,
x"02" after 7670950 ns,
x"23" after 7681800 ns,
x"88" after 7692650 ns,
x"E7" after 7703500 ns,
x"FC" after 7714350 ns,
x"83" after 7725200 ns,
x"27" after 7736050 ns,
x"44" after 7746900 ns,
x"FF" after 7757750 ns,
x"23" after 7768600 ns,
x"26" after 7779450 ns,
x"F4" after 7790300 ns,
x"FE" after 7801150 ns,
x"23" after 7812000 ns,
x"28" after 7822850 ns,
x"04" after 7833700 ns,
x"FE" after 7844550 ns,
x"6F" after 7855400 ns,
x"00" after 7866250 ns,
x"C0" after 7877100 ns,
x"03" after 7887950 ns,
x"83" after 7898800 ns,
x"27" after 7909650 ns,
x"C4" after 7920500 ns,
x"FE" after 7931350 ns,
x"13" after 7942200 ns,
x"87" after 7953050 ns,
x"F7" after 7963900 ns,
x"FF" after 7974750 ns,
x"83" after 7985600 ns,
x"27" after 7996450 ns,
x"04" after 8007300 ns,
x"FF" after 8018150 ns,
x"33" after 8029000 ns,
x"07" after 8039850 ns,
x"F7" after 8050700 ns,
x"40" after 8061550 ns,
x"83" after 8072400 ns,
x"27" after 8083250 ns,
x"04" after 8094100 ns,
x"FF" after 8104950 ns,
x"83" after 8115800 ns,
x"26" after 8126650 ns,
x"44" after 8137500 ns,
x"FC" after 8148350 ns,
x"B3" after 8159200 ns,
x"87" after 8170050 ns,
x"F6" after 8180900 ns,
x"00" after 8191750 ns,
x"13" after 8202600 ns,
x"07" after 8213450 ns,
x"87" after 8224300 ns,
x"FF" after 8235150 ns,
x"33" after 8246000 ns,
x"07" after 8256850 ns,
x"87" after 8267700 ns,
x"00" after 8278550 ns,
x"03" after 8289400 ns,
x"47" after 8300250 ns,
x"07" after 8311100 ns,
x"FD" after 8321950 ns,
x"23" after 8332800 ns,
x"80" after 8343650 ns,
x"E7" after 8354500 ns,
x"00" after 8365350 ns,
x"83" after 8376200 ns,
x"27" after 8387050 ns,
x"04" after 8397900 ns,
x"FF" after 8408750 ns,
x"93" after 8419600 ns,
x"87" after 8430450 ns,
x"17" after 8441300 ns,
x"00" after 8452150 ns,
x"23" after 8463000 ns,
x"28" after 8473850 ns,
x"F4" after 8484700 ns,
x"FE" after 8495550 ns,
x"03" after 8506400 ns,
x"27" after 8517250 ns,
x"04" after 8528100 ns,
x"FF" after 8538950 ns,
x"83" after 8549800 ns,
x"27" after 8560650 ns,
x"C4" after 8571500 ns,
x"FE" after 8582350 ns,
x"E3" after 8593200 ns,
x"40" after 8604050 ns,
x"F7" after 8614900 ns,
x"FC" after 8625750 ns,
x"83" after 8636600 ns,
x"27" after 8647450 ns,
x"C4" after 8658300 ns,
x"FE" after 8669150 ns,
x"03" after 8680000 ns,
x"27" after 8690850 ns,
x"44" after 8701700 ns,
x"FC" after 8712550 ns,
x"B3" after 8723400 ns,
x"07" after 8734250 ns,
x"F7" after 8745100 ns,
x"00" after 8755950 ns,
x"23" after 8766800 ns,
x"80" after 8777650 ns,
x"07" after 8788500 ns,
x"00" after 8799350 ns,
x"83" after 8810200 ns,
x"27" after 8821050 ns,
x"C4" after 8831900 ns,
x"FE" after 8842750 ns,
x"13" after 8853600 ns,
x"85" after 8864450 ns,
x"07" after 8875300 ns,
x"00" after 8886150 ns,
x"03" after 8897000 ns,
x"24" after 8907850 ns,
x"C1" after 8918700 ns,
x"03" after 8929550 ns,
x"13" after 8940400 ns,
x"01" after 8951250 ns,
x"01" after 8962100 ns,
x"04" after 8972950 ns,
x"67" after 8983800 ns,
x"80" after 8994650 ns,
x"00" after 9005500 ns,
x"00" after 9016350 ns,
x"13" after 9027200 ns,
x"01" after 9038050 ns,
x"01" after 9048900 ns,
x"FB" after 9059750 ns,
x"23" after 9070600 ns,
x"2A" after 9081450 ns,
x"11" after 9092300 ns,
x"02" after 9103150 ns,
x"23" after 9114000 ns,
x"28" after 9124850 ns,
x"81" after 9135700 ns,
x"02" after 9146550 ns,
x"13" after 9157400 ns,
x"04" after 9168250 ns,
x"81" after 9179100 ns,
x"03" after 9189950 ns,
x"23" after 9200800 ns,
x"2A" after 9211650 ns,
x"A4" after 9222500 ns,
x"FC" after 9233350 ns,
x"23" after 9244200 ns,
x"28" after 9255050 ns,
x"B4" after 9265900 ns,
x"FC" after 9276750 ns,
x"23" after 9287600 ns,
x"20" after 9298450 ns,
x"C4" after 9309300 ns,
x"00" after 9320150 ns,
x"23" after 9331000 ns,
x"22" after 9341850 ns,
x"D4" after 9352700 ns,
x"00" after 9363550 ns,
x"23" after 9374400 ns,
x"24" after 9385250 ns,
x"E4" after 9396100 ns,
x"00" after 9406950 ns,
x"23" after 9417800 ns,
x"26" after 9428650 ns,
x"F4" after 9439500 ns,
x"00" after 9450350 ns,
x"23" after 9461200 ns,
x"28" after 9472050 ns,
x"04" after 9482900 ns,
x"01" after 9493750 ns,
x"23" after 9504600 ns,
x"2A" after 9515450 ns,
x"14" after 9526300 ns,
x"01" after 9537150 ns,
x"93" after 9548000 ns,
x"07" after 9558850 ns,
x"84" after 9569700 ns,
x"01" after 9580550 ns,
x"23" after 9591400 ns,
x"26" after 9602250 ns,
x"F4" after 9613100 ns,
x"FC" after 9623950 ns,
x"83" after 9634800 ns,
x"27" after 9645650 ns,
x"C4" after 9656500 ns,
x"FC" after 9667350 ns,
x"93" after 9678200 ns,
x"87" after 9689050 ns,
x"87" after 9699900 ns,
x"FE" after 9710750 ns,
x"23" after 9721600 ns,
x"2E" after 9732450 ns,
x"F4" after 9743300 ns,
x"FC" after 9754150 ns,
x"83" after 9765000 ns,
x"27" after 9775850 ns,
x"04" after 9786700 ns,
x"FD" after 9797550 ns,
x"23" after 9808400 ns,
x"2A" after 9819250 ns,
x"F4" after 9830100 ns,
x"FE" after 9840950 ns,
x"83" after 9851800 ns,
x"27" after 9862650 ns,
x"44" after 9873500 ns,
x"FD" after 9884350 ns,
x"23" after 9895200 ns,
x"28" after 9906050 ns,
x"F4" after 9916900 ns,
x"FE" after 9927750 ns,
x"6F" after 9938600 ns,
x"00" after 9949450 ns,
x"00" after 9960300 ns,
x"21" after 9971150 ns,
x"83" after 9982000 ns,
x"27" after 9992850 ns,
x"44" after 10003700 ns,
x"FF" after 10014550 ns,
x"03" after 10025400 ns,
x"C7" after 10036250 ns,
x"07" after 10047100 ns,
x"00" after 10057950 ns,
x"93" after 10068800 ns,
x"07" after 10079650 ns,
x"50" after 10090500 ns,
x"02" after 10101350 ns,
x"63" after 10112200 ns,
x"1E" after 10123050 ns,
x"F7" after 10133900 ns,
x"1C" after 10144750 ns,
x"83" after 10155600 ns,
x"27" after 10166450 ns,
x"44" after 10177300 ns,
x"FF" after 10188150 ns,
x"93" after 10199000 ns,
x"87" after 10209850 ns,
x"17" after 10220700 ns,
x"00" after 10231550 ns,
x"23" after 10242400 ns,
x"2A" after 10253250 ns,
x"F4" after 10264100 ns,
x"FE" after 10274950 ns,
x"83" after 10285800 ns,
x"27" after 10296650 ns,
x"44" after 10307500 ns,
x"FF" after 10318350 ns,
x"83" after 10329200 ns,
x"C7" after 10340050 ns,
x"07" after 10350900 ns,
x"00" after 10361750 ns,
x"13" after 10372600 ns,
x"07" after 10383450 ns,
x"30" after 10394300 ns,
x"07" after 10405150 ns,
x"63" after 10416000 ns,
x"8C" after 10426850 ns,
x"E7" after 10437700 ns,
x"06" after 10448550 ns,
x"13" after 10459400 ns,
x"07" after 10470250 ns,
x"30" after 10481100 ns,
x"07" after 10491950 ns,
x"63" after 10502800 ns,
x"44" after 10513650 ns,
x"F7" after 10524500 ns,
x"18" after 10535350 ns,
x"13" after 10546200 ns,
x"07" after 10557050 ns,
x"40" after 10567900 ns,
x"06" after 10578750 ns,
x"63" after 10589600 ns,
x"88" after 10600450 ns,
x"E7" after 10611300 ns,
x"02" after 10622150 ns,
x"13" after 10633000 ns,
x"07" after 10643850 ns,
x"40" after 10654700 ns,
x"06" after 10665550 ns,
x"63" after 10676400 ns,
x"4C" after 10687250 ns,
x"F7" after 10698100 ns,
x"16" after 10708950 ns,
x"13" after 10719800 ns,
x"07" after 10730650 ns,
x"30" after 10741500 ns,
x"06" after 10752350 ns,
x"63" after 10763200 ns,
x"88" after 10774050 ns,
x"E7" after 10784900 ns,
x"08" after 10795750 ns,
x"13" after 10806600 ns,
x"07" after 10817450 ns,
x"30" after 10828300 ns,
x"06" after 10839150 ns,
x"63" after 10850000 ns,
x"44" after 10860850 ns,
x"F7" after 10871700 ns,
x"16" after 10882550 ns,
x"13" after 10893400 ns,
x"07" after 10904250 ns,
x"50" after 10915100 ns,
x"02" after 10925950 ns,
x"63" after 10936800 ns,
x"86" after 10947650 ns,
x"E7" after 10958500 ns,
x"0A" after 10969350 ns,
x"13" after 10980200 ns,
x"07" after 10991050 ns,
x"00" after 11001900 ns,
x"03" after 11012750 ns,
x"63" after 11023600 ns,
x"8E" after 11034450 ns,
x"E7" after 11045300 ns,
x"0A" after 11056150 ns,
x"6F" after 11067000 ns,
x"00" after 11077850 ns,
x"40" after 11088700 ns,
x"15" after 11099550 ns,
x"83" after 11110400 ns,
x"27" after 11121250 ns,
x"C4" after 11132100 ns,
x"FD" after 11142950 ns,
x"13" after 11153800 ns,
x"87" after 11164650 ns,
x"47" after 11175500 ns,
x"00" after 11186350 ns,
x"23" after 11197200 ns,
x"2E" after 11208050 ns,
x"E4" after 11218900 ns,
x"FC" after 11229750 ns,
x"83" after 11240600 ns,
x"A7" after 11251450 ns,
x"07" after 11262300 ns,
x"00" after 11273150 ns,
x"23" after 11284000 ns,
x"24" after 11294850 ns,
x"F4" after 11305700 ns,
x"FE" after 11316550 ns,
x"83" after 11327400 ns,
x"25" after 11338250 ns,
x"84" after 11349100 ns,
x"FE" after 11359950 ns,
x"03" after 11370800 ns,
x"25" after 11381650 ns,
x"04" after 11392500 ns,
x"FF" after 11403350 ns,
x"EF" after 11414200 ns,
x"F0" after 11425050 ns,
x"1F" after 11435900 ns,
x"E0" after 11446750 ns,
x"93" after 11457600 ns,
x"07" after 11468450 ns,
x"05" after 11479300 ns,
x"00" after 11490150 ns,
x"13" after 11501000 ns,
x"87" after 11511850 ns,
x"07" after 11522700 ns,
x"00" after 11533550 ns,
x"83" after 11544400 ns,
x"27" after 11555250 ns,
x"04" after 11566100 ns,
x"FF" after 11576950 ns,
x"B3" after 11587800 ns,
x"87" after 11598650 ns,
x"E7" after 11609500 ns,
x"00" after 11620350 ns,
x"23" after 11631200 ns,
x"28" after 11642050 ns,
x"F4" after 11652900 ns,
x"FE" after 11663750 ns,
x"6F" after 11674600 ns,
x"00" after 11685450 ns,
x"40" after 11696300 ns,
x"16" after 11707150 ns,
x"83" after 11718000 ns,
x"27" after 11728850 ns,
x"C4" after 11739700 ns,
x"FD" after 11750550 ns,
x"13" after 11761400 ns,
x"87" after 11772250 ns,
x"47" after 11783100 ns,
x"00" after 11793950 ns,
x"23" after 11804800 ns,
x"2E" after 11815650 ns,
x"E4" after 11826500 ns,
x"FC" after 11837350 ns,
x"83" after 11848200 ns,
x"A7" after 11859050 ns,
x"07" after 11869900 ns,
x"00" after 11880750 ns,
x"23" after 11891600 ns,
x"26" after 11902450 ns,
x"F4" after 11913300 ns,
x"FE" after 11924150 ns,
x"83" after 11935000 ns,
x"25" after 11945850 ns,
x"C4" after 11956700 ns,
x"FE" after 11967550 ns,
x"03" after 11978400 ns,
x"25" after 11989250 ns,
x"04" after 12000100 ns,
x"FF" after 12010950 ns,
x"EF" after 12021800 ns,
x"F0" after 12032650 ns,
x"5F" after 12043500 ns,
x"CB" after 12054350 ns,
x"93" after 12065200 ns,
x"07" after 12076050 ns,
x"05" after 12086900 ns,
x"00" after 12097750 ns,
x"13" after 12108600 ns,
x"87" after 12119450 ns,
x"07" after 12130300 ns,
x"00" after 12141150 ns,
x"83" after 12152000 ns,
x"27" after 12162850 ns,
x"04" after 12173700 ns,
x"FF" after 12184550 ns,
x"B3" after 12195400 ns,
x"87" after 12206250 ns,
x"E7" after 12217100 ns,
x"00" after 12227950 ns,
x"23" after 12238800 ns,
x"28" after 12249650 ns,
x"F4" after 12260500 ns,
x"FE" after 12271350 ns,
x"6F" after 12282200 ns,
x"00" after 12293050 ns,
x"C0" after 12303900 ns,
x"12" after 12314750 ns,
x"83" after 12325600 ns,
x"27" after 12336450 ns,
x"C4" after 12347300 ns,
x"FD" after 12358150 ns,
x"13" after 12369000 ns,
x"87" after 12379850 ns,
x"47" after 12390700 ns,
x"00" after 12401550 ns,
x"23" after 12412400 ns,
x"2E" after 12423250 ns,
x"E4" after 12434100 ns,
x"FC" after 12444950 ns,
x"83" after 12455800 ns,
x"A7" after 12466650 ns,
x"07" after 12477500 ns,
x"00" after 12488350 ns,
x"A3" after 12499200 ns,
x"03" after 12510050 ns,
x"F4" after 12520900 ns,
x"FE" after 12531750 ns,
x"83" after 12542600 ns,
x"27" after 12553450 ns,
x"04" after 12564300 ns,
x"FF" after 12575150 ns,
x"13" after 12586000 ns,
x"87" after 12596850 ns,
x"17" after 12607700 ns,
x"00" after 12618550 ns,
x"23" after 12629400 ns,
x"28" after 12640250 ns,
x"E4" after 12651100 ns,
x"FE" after 12661950 ns,
x"03" after 12672800 ns,
x"47" after 12683650 ns,
x"74" after 12694500 ns,
x"FE" after 12705350 ns,
x"23" after 12716200 ns,
x"80" after 12727050 ns,
x"E7" after 12737900 ns,
x"00" after 12748750 ns,
x"6F" after 12759600 ns,
x"00" after 12770450 ns,
x"00" after 12781300 ns,
x"10" after 12792150 ns,
x"83" after 12803000 ns,
x"27" after 12813850 ns,
x"04" after 12824700 ns,
x"FF" after 12835550 ns,
x"13" after 12846400 ns,
x"87" after 12857250 ns,
x"17" after 12868100 ns,
x"00" after 12878950 ns,
x"23" after 12889800 ns,
x"28" after 12900650 ns,
x"E4" after 12911500 ns,
x"FE" after 12922350 ns,
x"13" after 12933200 ns,
x"07" after 12944050 ns,
x"50" after 12954900 ns,
x"02" after 12965750 ns,
x"23" after 12976600 ns,
x"80" after 12987450 ns,
x"E7" after 12998300 ns,
x"00" after 13009150 ns,
x"6F" after 13020000 ns,
x"00" after 13030850 ns,
x"80" after 13041700 ns,
x"0E" after 13052550 ns,
x"83" after 13063400 ns,
x"27" after 13074250 ns,
x"44" after 13085100 ns,
x"FF" after 13095950 ns,
x"93" after 13106800 ns,
x"87" after 13117650 ns,
x"17" after 13128500 ns,
x"00" after 13139350 ns,
x"03" after 13150200 ns,
x"C7" after 13161050 ns,
x"07" after 13171900 ns,
x"00" after 13182750 ns,
x"93" after 13193600 ns,
x"07" after 13204450 ns,
x"20" after 13215300 ns,
x"03" after 13226150 ns,
x"63" after 13237000 ns,
x"10" after 13247850 ns,
x"F7" after 13258700 ns,
x"06" after 13269550 ns,
x"83" after 13280400 ns,
x"27" after 13291250 ns,
x"44" after 13302100 ns,
x"FF" after 13312950 ns,
x"93" after 13323800 ns,
x"87" after 13334650 ns,
x"27" after 13345500 ns,
x"00" after 13356350 ns,
x"03" after 13367200 ns,
x"C7" after 13378050 ns,
x"07" after 13388900 ns,
x"00" after 13399750 ns,
x"93" after 13410600 ns,
x"07" after 13421450 ns,
x"80" after 13432300 ns,
x"05" after 13443150 ns,
x"63" after 13454000 ns,
x"16" after 13464850 ns,
x"F7" after 13475700 ns,
x"04" after 13486550 ns,
x"83" after 13497400 ns,
x"27" after 13508250 ns,
x"44" after 13519100 ns,
x"FF" after 13529950 ns,
x"93" after 13540800 ns,
x"87" after 13551650 ns,
x"27" after 13562500 ns,
x"00" after 13573350 ns,
x"23" after 13584200 ns,
x"2A" after 13595050 ns,
x"F4" after 13605900 ns,
x"FE" after 13616750 ns,
x"83" after 13627600 ns,
x"27" after 13638450 ns,
x"C4" after 13649300 ns,
x"FD" after 13660150 ns,
x"13" after 13671000 ns,
x"87" after 13681850 ns,
x"47" after 13692700 ns,
x"00" after 13703550 ns,
x"23" after 13714400 ns,
x"2E" after 13725250 ns,
x"E4" after 13736100 ns,
x"FC" after 13746950 ns,
x"83" after 13757800 ns,
x"A7" after 13768650 ns,
x"07" after 13779500 ns,
x"00" after 13790350 ns,
x"23" after 13801200 ns,
x"20" after 13812050 ns,
x"F4" after 13822900 ns,
x"FE" after 13833750 ns,
x"83" after 13844600 ns,
x"25" after 13855450 ns,
x"04" after 13866300 ns,
x"FE" after 13877150 ns,
x"03" after 13888000 ns,
x"25" after 13898850 ns,
x"04" after 13909700 ns,
x"FF" after 13920550 ns,
x"EF" after 13931400 ns,
x"F0" after 13942250 ns,
x"5F" after 13953100 ns,
x"C7" after 13963950 ns,
x"93" after 13974800 ns,
x"07" after 13985650 ns,
x"05" after 13996500 ns,
x"00" after 14007350 ns,
x"13" after 14018200 ns,
x"87" after 14029050 ns,
x"07" after 14039900 ns,
x"00" after 14050750 ns,
x"83" after 14061600 ns,
x"27" after 14072450 ns,
x"04" after 14083300 ns,
x"FF" after 14094150 ns,
x"B3" after 14105000 ns,
x"87" after 14115850 ns,
x"E7" after 14126700 ns,
x"00" after 14137550 ns,
x"23" after 14148400 ns,
x"28" after 14159250 ns,
x"F4" after 14170100 ns,
x"FE" after 14180950 ns,
x"13" after 14191800 ns,
x"00" after 14202650 ns,
x"00" after 14213500 ns,
x"00" after 14224350 ns,
x"6F" after 14235200 ns,
x"00" after 14246050 ns,
x"80" after 14256900 ns,
x"07" after 14267750 ns,
x"83" after 14278600 ns,
x"27" after 14289450 ns,
x"04" after 14300300 ns,
x"FF" after 14311150 ns,
x"13" after 14322000 ns,
x"87" after 14332850 ns,
x"17" after 14343700 ns,
x"00" after 14354550 ns,
x"23" after 14365400 ns,
x"28" after 14376250 ns,
x"E4" after 14387100 ns,
x"FE" after 14397950 ns,
x"13" after 14408800 ns,
x"07" after 14419650 ns,
x"50" after 14430500 ns,
x"02" after 14441350 ns,
x"23" after 14452200 ns,
x"80" after 14463050 ns,
x"E7" after 14473900 ns,
x"00" after 14484750 ns,
x"83" after 14495600 ns,
x"27" after 14506450 ns,
x"04" after 14517300 ns,
x"FF" after 14528150 ns,
x"13" after 14539000 ns,
x"87" after 14549850 ns,
x"17" after 14560700 ns,
x"00" after 14571550 ns,
x"23" after 14582400 ns,
x"28" after 14593250 ns,
x"E4" after 14604100 ns,
x"FE" after 14614950 ns,
x"13" after 14625800 ns,
x"07" after 14636650 ns,
x"00" after 14647500 ns,
x"03" after 14658350 ns,
x"23" after 14669200 ns,
x"80" after 14680050 ns,
x"E7" after 14690900 ns,
x"00" after 14701750 ns,
x"6F" after 14712600 ns,
x"00" after 14723450 ns,
x"C0" after 14734300 ns,
x"04" after 14745150 ns,
x"83" after 14756000 ns,
x"27" after 14766850 ns,
x"04" after 14777700 ns,
x"FF" after 14788550 ns,
x"13" after 14799400 ns,
x"87" after 14810250 ns,
x"17" after 14821100 ns,
x"00" after 14831950 ns,
x"23" after 14842800 ns,
x"28" after 14853650 ns,
x"E4" after 14864500 ns,
x"FE" after 14875350 ns,
x"13" after 14886200 ns,
x"07" after 14897050 ns,
x"50" after 14907900 ns,
x"02" after 14918750 ns,
x"23" after 14929600 ns,
x"80" after 14940450 ns,
x"E7" after 14951300 ns,
x"00" after 14962150 ns,
x"83" after 14973000 ns,
x"27" after 14983850 ns,
x"04" after 14994700 ns,
x"FF" after 15005550 ns,
x"13" after 15016400 ns,
x"87" after 15027250 ns,
x"17" after 15038100 ns,
x"00" after 15048950 ns,
x"23" after 15059800 ns,
x"28" after 15070650 ns,
x"E4" after 15081500 ns,
x"FE" after 15092350 ns,
x"03" after 15103200 ns,
x"27" after 15114050 ns,
x"44" after 15124900 ns,
x"FF" after 15135750 ns,
x"03" after 15146600 ns,
x"47" after 15157450 ns,
x"07" after 15168300 ns,
x"00" after 15179150 ns,
x"23" after 15190000 ns,
x"80" after 15200850 ns,
x"E7" after 15211700 ns,
x"00" after 15222550 ns,
x"6F" after 15233400 ns,
x"00" after 15244250 ns,
x"C0" after 15255100 ns,
x"01" after 15265950 ns,
x"83" after 15276800 ns,
x"27" after 15287650 ns,
x"04" after 15298500 ns,
x"FF" after 15309350 ns,
x"13" after 15320200 ns,
x"87" after 15331050 ns,
x"17" after 15341900 ns,
x"00" after 15352750 ns,
x"23" after 15363600 ns,
x"28" after 15374450 ns,
x"E4" after 15385300 ns,
x"FE" after 15396150 ns,
x"03" after 15407000 ns,
x"27" after 15417850 ns,
x"44" after 15428700 ns,
x"FF" after 15439550 ns,
x"03" after 15450400 ns,
x"47" after 15461250 ns,
x"07" after 15472100 ns,
x"00" after 15482950 ns,
x"23" after 15493800 ns,
x"80" after 15504650 ns,
x"E7" after 15515500 ns,
x"00" after 15526350 ns,
x"83" after 15537200 ns,
x"27" after 15548050 ns,
x"44" after 15558900 ns,
x"FF" after 15569750 ns,
x"93" after 15580600 ns,
x"87" after 15591450 ns,
x"17" after 15602300 ns,
x"00" after 15613150 ns,
x"23" after 15624000 ns,
x"2A" after 15634850 ns,
x"F4" after 15645700 ns,
x"FE" after 15656550 ns,
x"83" after 15667400 ns,
x"27" after 15678250 ns,
x"44" after 15689100 ns,
x"FF" after 15699950 ns,
x"83" after 15710800 ns,
x"C7" after 15721650 ns,
x"07" after 15732500 ns,
x"00" after 15743350 ns,
x"E3" after 15754200 ns,
x"96" after 15765050 ns,
x"07" after 15775900 ns,
x"DE" after 15786750 ns,
x"83" after 15797600 ns,
x"27" after 15808450 ns,
x"04" after 15819300 ns,
x"FF" after 15830150 ns,
x"23" after 15841000 ns,
x"80" after 15851850 ns,
x"07" after 15862700 ns,
x"00" after 15873550 ns,
x"13" after 15884400 ns,
x"00" after 15895250 ns,
x"00" after 15906100 ns,
x"00" after 15916950 ns,
x"83" after 15927800 ns,
x"20" after 15938650 ns,
x"41" after 15949500 ns,
x"03" after 15960350 ns,
x"03" after 15971200 ns,
x"24" after 15982050 ns,
x"01" after 15992900 ns,
x"03" after 16003750 ns,
x"13" after 16014600 ns,
x"01" after 16025450 ns,
x"01" after 16036300 ns,
x"05" after 16047150 ns,
x"67" after 16058000 ns,
x"80" after 16068850 ns,
x"00" after 16079700 ns,
x"00" after 16090550 ns,
x"13" after 16101400 ns,
x"01" after 16112250 ns,
x"01" after 16123100 ns,
x"FF" after 16133950 ns,
x"23" after 16144800 ns,
x"26" after 16155650 ns,
x"11" after 16166500 ns,
x"00" after 16177350 ns,
x"23" after 16188200 ns,
x"24" after 16199050 ns,
x"81" after 16209900 ns,
x"00" after 16220750 ns,
x"13" after 16231600 ns,
x"04" after 16242450 ns,
x"01" after 16253300 ns,
x"01" after 16264150 ns,
x"13" after 16275000 ns,
x"05" after 16285850 ns,
x"00" after 16296700 ns,
x"00" after 16307550 ns,
x"EF" after 16318400 ns,
x"F0" after 16329250 ns,
x"DF" after 16340100 ns,
x"AC" after 16350950 ns,
x"93" after 16361800 ns,
x"07" after 16372650 ns,
x"05" after 16383500 ns,
x"00" after 16394350 ns,
x"A3" after 16405200 ns,
x"0B" after 16416050 ns,
x"F4" after 16426900 ns,
x"FE" after 16437750 ns,
x"03" after 16448600 ns,
x"47" after 16459450 ns,
x"74" after 16470300 ns,
x"FF" after 16481150 ns,
x"93" after 16492000 ns,
x"07" after 16502850 ns,
x"D0" after 16513700 ns,
x"00" after 16524550 ns,
x"63" after 16535400 ns,
x"1E" after 16546250 ns,
x"F7" after 16557100 ns,
x"04" after 16567950 ns,
x"B7" after 16578800 ns,
x"17" after 16589650 ns,
x"00" after 16600500 ns,
x"00" after 16611350 ns,
x"83" after 16622200 ns,
x"A7" after 16633050 ns,
x"07" after 16643900 ns,
x"80" after 16654750 ns,
x"93" after 16665600 ns,
x"86" after 16676450 ns,
x"17" after 16687300 ns,
x"00" after 16698150 ns,
x"37" after 16709000 ns,
x"17" after 16719850 ns,
x"00" after 16730700 ns,
x"00" after 16741550 ns,
x"23" after 16752400 ns,
x"20" after 16763250 ns,
x"D7" after 16774100 ns,
x"80" after 16784950 ns,
x"37" after 16795800 ns,
x"17" after 16806650 ns,
x"00" after 16817500 ns,
x"00" after 16828350 ns,
x"13" after 16839200 ns,
x"07" after 16850050 ns,
x"47" after 16860900 ns,
x"8C" after 16871750 ns,
x"B3" after 16882600 ns,
x"07" after 16893450 ns,
x"F7" after 16904300 ns,
x"00" after 16915150 ns,
x"03" after 16926000 ns,
x"47" after 16936850 ns,
x"74" after 16947700 ns,
x"FF" after 16958550 ns,
x"23" after 16969400 ns,
x"80" after 16980250 ns,
x"E7" after 16991100 ns,
x"00" after 17001950 ns,
x"B7" after 17012800 ns,
x"17" after 17023650 ns,
x"00" after 17034500 ns,
x"00" after 17045350 ns,
x"83" after 17056200 ns,
x"A7" after 17067050 ns,
x"07" after 17077900 ns,
x"80" after 17088750 ns,
x"93" after 17099600 ns,
x"86" after 17110450 ns,
x"17" after 17121300 ns,
x"00" after 17132150 ns,
x"37" after 17143000 ns,
x"17" after 17153850 ns,
x"00" after 17164700 ns,
x"00" after 17175550 ns,
x"23" after 17186400 ns,
x"20" after 17197250 ns,
x"D7" after 17208100 ns,
x"80" after 17218950 ns,
x"37" after 17229800 ns,
x"17" after 17240650 ns,
x"00" after 17251500 ns,
x"00" after 17262350 ns,
x"13" after 17273200 ns,
x"07" after 17284050 ns,
x"47" after 17294900 ns,
x"8C" after 17305750 ns,
x"B3" after 17316600 ns,
x"07" after 17327450 ns,
x"F7" after 17338300 ns,
x"00" after 17349150 ns,
x"23" after 17360000 ns,
x"80" after 17370850 ns,
x"07" after 17381700 ns,
x"00" after 17392550 ns,
x"B7" after 17403400 ns,
x"17" after 17414250 ns,
x"00" after 17425100 ns,
x"00" after 17435950 ns,
x"13" after 17446800 ns,
x"07" after 17457650 ns,
x"10" after 17468500 ns,
x"00" after 17479350 ns,
x"23" after 17490200 ns,
x"A2" after 17501050 ns,
x"E7" after 17511900 ns,
x"80" after 17522750 ns,
x"B7" after 17533600 ns,
x"17" after 17544450 ns,
x"00" after 17555300 ns,
x"00" after 17566150 ns,
x"83" after 17577000 ns,
x"A7" after 17587850 ns,
x"07" after 17598700 ns,
x"80" after 17609550 ns,
x"93" after 17620400 ns,
x"86" after 17631250 ns,
x"17" after 17642100 ns,
x"00" after 17652950 ns,
x"37" after 17663800 ns,
x"17" after 17674650 ns,
x"00" after 17685500 ns,
x"00" after 17696350 ns,
x"23" after 17707200 ns,
x"20" after 17718050 ns,
x"D7" after 17728900 ns,
x"80" after 17739750 ns,
x"37" after 17750600 ns,
x"17" after 17761450 ns,
x"00" after 17772300 ns,
x"00" after 17783150 ns,
x"13" after 17794000 ns,
x"07" after 17804850 ns,
x"47" after 17815700 ns,
x"8C" after 17826550 ns,
x"B3" after 17837400 ns,
x"07" after 17848250 ns,
x"F7" after 17859100 ns,
x"00" after 17869950 ns,
x"03" after 17880800 ns,
x"47" after 17891650 ns,
x"74" after 17902500 ns,
x"FF" after 17913350 ns,
x"23" after 17924200 ns,
x"80" after 17935050 ns,
x"E7" after 17945900 ns,
x"00" after 17956750 ns,
x"13" after 17967600 ns,
x"00" after 17978450 ns,
x"00" after 17989300 ns,
x"00" after 18000150 ns,
x"83" after 18011000 ns,
x"20" after 18021850 ns,
x"C1" after 18032700 ns,
x"00" after 18043550 ns,
x"03" after 18054400 ns,
x"24" after 18065250 ns,
x"81" after 18076100 ns,
x"00" after 18086950 ns,
x"13" after 18097800 ns,
x"01" after 18108650 ns,
x"01" after 18119500 ns,
x"01" after 18130350 ns,
x"67" after 18141200 ns,
x"80" after 18152050 ns,
x"00" after 18162900 ns,
x"00" after 18173750 ns,
x"13" after 18184600 ns,
x"01" after 18195450 ns,
x"81" after 18206300 ns,
x"FE" after 18217150 ns,
x"23" after 18228000 ns,
x"2A" after 18238850 ns,
x"81" after 18249700 ns,
x"00" after 18260550 ns,
x"13" after 18271400 ns,
x"04" after 18282250 ns,
x"81" after 18293100 ns,
x"01" after 18303950 ns,
x"23" after 18314800 ns,
x"26" after 18325650 ns,
x"A4" after 18336500 ns,
x"FE" after 18347350 ns,
x"B7" after 18358200 ns,
x"17" after 18369050 ns,
x"00" after 18379900 ns,
x"00" after 18390750 ns,
x"83" after 18401600 ns,
x"A7" after 18412450 ns,
x"47" after 18423300 ns,
x"80" after 18434150 ns,
x"63" after 18445000 ns,
x"96" after 18455850 ns,
x"07" after 18466700 ns,
x"00" after 18477550 ns,
x"93" after 18488400 ns,
x"07" after 18499250 ns,
x"00" after 18510100 ns,
x"00" after 18520950 ns,
x"6F" after 18531800 ns,
x"00" after 18542650 ns,
x"40" after 18553500 ns,
x"03" after 18564350 ns,
x"83" after 18575200 ns,
x"27" after 18586050 ns,
x"C4" after 18596900 ns,
x"FE" after 18607750 ns,
x"37" after 18618600 ns,
x"17" after 18629450 ns,
x"00" after 18640300 ns,
x"00" after 18651150 ns,
x"13" after 18662000 ns,
x"07" after 18672850 ns,
x"47" after 18683700 ns,
x"8C" after 18694550 ns,
x"23" after 18705400 ns,
x"A0" after 18716250 ns,
x"E7" after 18727100 ns,
x"00" after 18737950 ns,
x"B7" after 18748800 ns,
x"17" after 18759650 ns,
x"00" after 18770500 ns,
x"00" after 18781350 ns,
x"83" after 18792200 ns,
x"A7" after 18803050 ns,
x"07" after 18813900 ns,
x"80" after 18824750 ns,
x"23" after 18835600 ns,
x"2A" after 18846450 ns,
x"F4" after 18857300 ns,
x"FE" after 18868150 ns,
x"B7" after 18879000 ns,
x"17" after 18889850 ns,
x"00" after 18900700 ns,
x"00" after 18911550 ns,
x"23" after 18922400 ns,
x"A0" after 18933250 ns,
x"07" after 18944100 ns,
x"80" after 18954950 ns,
x"B7" after 18965800 ns,
x"17" after 18976650 ns,
x"00" after 18987500 ns,
x"00" after 18998350 ns,
x"23" after 19009200 ns,
x"A2" after 19020050 ns,
x"07" after 19030900 ns,
x"80" after 19041750 ns,
x"83" after 19052600 ns,
x"27" after 19063450 ns,
x"44" after 19074300 ns,
x"FF" after 19085150 ns,
x"13" after 19096000 ns,
x"85" after 19106850 ns,
x"07" after 19117700 ns,
x"00" after 19128550 ns,
x"03" after 19139400 ns,
x"24" after 19150250 ns,
x"41" after 19161100 ns,
x"01" after 19171950 ns,
x"13" after 19182800 ns,
x"01" after 19193650 ns,
x"81" after 19204500 ns,
x"01" after 19215350 ns,
x"67" after 19226200 ns,
x"80" after 19237050 ns,
x"00" after 19247900 ns,
x"00" after 19258750 ns,
x"13" after 19269600 ns,
x"01" after 19280450 ns,
x"01" after 19291300 ns,
x"FF" after 19302150 ns,
x"23" after 19313000 ns,
x"26" after 19323850 ns,
x"11" after 19334700 ns,
x"00" after 19345550 ns,
x"23" after 19356400 ns,
x"24" after 19367250 ns,
x"81" after 19378100 ns,
x"00" after 19388950 ns,
x"13" after 19399800 ns,
x"04" after 19410650 ns,
x"01" after 19421500 ns,
x"01" after 19432350 ns,
x"B7" after 19443200 ns,
x"27" after 19454050 ns,
x"00" after 19464900 ns,
x"00" after 19475750 ns,
x"93" after 19486600 ns,
x"85" after 19497450 ns,
x"07" after 19508300 ns,
x"06" after 19519150 ns,
x"13" after 19530000 ns,
x"05" after 19540850 ns,
x"00" after 19551700 ns,
x"00" after 19562550 ns,
x"EF" after 19573400 ns,
x"F0" after 19584250 ns,
x"5F" after 19595100 ns,
x"93" after 19605950 ns,
x"B7" after 19616800 ns,
x"17" after 19627650 ns,
x"00" after 19638500 ns,
x"00" after 19649350 ns,
x"13" after 19660200 ns,
x"85" after 19671050 ns,
x"C7" after 19681900 ns,
x"81" after 19692750 ns,
x"EF" after 19703600 ns,
x"F0" after 19714450 ns,
x"9F" after 19725300 ns,
x"98" after 19736150 ns,
x"13" after 19747000 ns,
x"05" after 19757850 ns,
x"10" after 19768700 ns,
x"00" after 19779550 ns,
x"EF" after 19790400 ns,
x"F0" after 19801250 ns,
x"5F" after 19812100 ns,
x"97" after 19822950 ns,
x"B7" after 19833800 ns,
x"17" after 19844650 ns,
x"00" after 19855500 ns,
x"00" after 19866350 ns,
x"13" after 19877200 ns,
x"85" after 19888050 ns,
x"47" after 19898900 ns,
x"83" after 19909750 ns,
x"EF" after 19920600 ns,
x"F0" after 19931450 ns,
x"5F" after 19942300 ns,
x"97" after 19953150 ns,
x"23" after 19964000 ns,
x"2A" after 19974850 ns,
x"04" after 19985700 ns,
x"FE" after 19996550 ns,
x"83" after 20007400 ns,
x"27" after 20018250 ns,
x"44" after 20029100 ns,
x"FF" after 20039950 ns,
x"93" after 20050800 ns,
x"87" after 20061650 ns,
x"17" after 20072500 ns,
x"00" after 20083350 ns,
x"23" after 20094200 ns,
x"2A" after 20105050 ns,
x"F4" after 20115900 ns,
x"FE" after 20126750 ns,
x"03" after 20137600 ns,
x"27" after 20148450 ns,
x"44" after 20159300 ns,
x"FF" after 20170150 ns,
x"93" after 20181000 ns,
x"07" after 20191850 ns,
x"50" after 20202700 ns,
x"00" after 20213550 ns,
x"E3" after 20224400 ns,
x"D6" after 20235250 ns,
x"E7" after 20246100 ns,
x"FE" after 20256950 ns,
x"23" after 20267800 ns,
x"28" after 20278650 ns,
x"04" after 20289500 ns,
x"FE" after 20300350 ns,
x"93" after 20311200 ns,
x"07" after 20322050 ns,
x"04" after 20332900 ns,
x"FF" after 20343750 ns,
x"13" after 20354600 ns,
x"85" after 20365450 ns,
x"07" after 20376300 ns,
x"00" after 20387150 ns,
x"EF" after 20398000 ns,
x"F0" after 20408850 ns,
x"5F" after 20419700 ns,
x"F3" after 20430550 ns,
x"93" after 20441400 ns,
x"07" after 20452250 ns,
x"05" after 20463100 ns,
x"00" after 20473950 ns,
x"E3" after 20484800 ns,
x"8A" after 20495650 ns,
x"07" after 20506500 ns,
x"FC" after 20517350 ns,
x"83" after 20528200 ns,
x"27" after 20539050 ns,
x"04" after 20549900 ns,
x"FF" after 20560750 ns,
x"13" after 20571600 ns,
x"85" after 20582450 ns,
x"07" after 20593300 ns,
x"00" after 20604150 ns,
x"EF" after 20615000 ns,
x"F0" after 20625850 ns,
x"5F" after 20636700 ns,
x"93" after 20647550 ns,
x"6F" after 20658400 ns,
x"F0" after 20669250 ns,
x"5F" after 20680100 ns,
x"FC" after 20690950 ns,
x"00" after 20701800 ns,
x"00" after 20712650 ns,
x"00" after 20723500 ns,
x"41" after 20734350 ns,
x"00" after 20745200 ns,
x"00" after 20756050 ns,
x"00" after 20766900 ns,
x"00" after 20777750 ns,
x"00" after 20788600 ns,
x"00" after 20799450 ns,
x"00" after 20810300 ns,
x"00" after 20821150 ns,
x"30" after 20832000 ns,
x"31" after 20842850 ns,
x"32" after 20853700 ns,
x"33" after 20864550 ns,
x"34" after 20875400 ns,
x"35" after 20886250 ns,
x"36" after 20897100 ns,
x"37" after 20907950 ns,
x"38" after 20918800 ns,
x"39" after 20929650 ns,
x"41" after 20940500 ns,
x"42" after 20951350 ns,
x"43" after 20962200 ns,
x"44" after 20973050 ns,
x"45" after 20983900 ns,
x"46" after 20994750 ns,
x"00" after 21005600 ns,
x"00" after 21016450 ns,
x"00" after 21027300 ns,
x"00" after 21038150 ns,
x"43" after 21049000 ns,
x"61" after 21059850 ns,
x"6C" after 21070700 ns,
x"6C" after 21081550 ns,
x"62" after 21092400 ns,
x"61" after 21103250 ns,
x"63" after 21114100 ns,
x"6B" after 21124950 ns,
x"20" after 21135800 ns,
x"72" after 21146650 ns,
x"65" after 21157500 ns,
x"67" after 21168350 ns,
x"69" after 21179200 ns,
x"73" after 21190050 ns,
x"74" after 21200900 ns,
x"65" after 21211750 ns,
x"72" after 21222600 ns,
x"65" after 21233450 ns,
x"64" after 21244300 ns,
x"20" after 21255150 ns,
x"0A" after 21266000 ns,
x"00" after 21276850 ns,
x"00" after 21287700 ns,
x"00" after 21298550 ns,
x"50" after 21309400 ns,
x"49" after 21320250 ns,
x"43" after 21331100 ns,
x"20" after 21341950 ns,
x"6D" after 21352800 ns,
x"61" after 21363650 ns,
x"73" after 21374500 ns,
x"6B" after 21385350 ns,
x"20" after 21396200 ns,
x"6F" after 21407050 ns,
x"6B" after 21417900 ns,
x"0A" after 21428750 ns,
x"00" after 21439600 ns, -- END OF PROGRAM
x"41" after 22201000 ns,
x"42" after 22213850 ns,
x"43" after 22224700 ns,
x"0D" after 22236550 ns;

-- VHDL for tx_dv:
tx_dv <= '1' after 0 ns, '0' after 50 ns,
'1' after 10850 ns, '0' after 10900 ns,
'1' after 21700 ns, '0' after 21750 ns,
'1' after 32550 ns, '0' after 32600 ns,
'1' after 43400 ns, '0' after 43450 ns,
'1' after 54250 ns, '0' after 54300 ns,
'1' after 65100 ns, '0' after 65150 ns,
'1' after 75950 ns, '0' after 76000 ns,
'1' after 86800 ns, '0' after 86850 ns,
'1' after 97650 ns, '0' after 97700 ns,
'1' after 108500 ns, '0' after 108550 ns,
'1' after 119350 ns, '0' after 119400 ns,
'1' after 130200 ns, '0' after 130250 ns,
'1' after 141050 ns, '0' after 141100 ns,
'1' after 151900 ns, '0' after 151950 ns,
'1' after 162750 ns, '0' after 162800 ns,
'1' after 173600 ns, '0' after 173650 ns,
'1' after 184450 ns, '0' after 184500 ns,
'1' after 195300 ns, '0' after 195350 ns,
'1' after 206150 ns, '0' after 206200 ns,
'1' after 217000 ns, '0' after 217050 ns,
'1' after 227850 ns, '0' after 227900 ns,
'1' after 238700 ns, '0' after 238750 ns,
'1' after 249550 ns, '0' after 249600 ns,
'1' after 260400 ns, '0' after 260450 ns,
'1' after 271250 ns, '0' after 271300 ns,
'1' after 282100 ns, '0' after 282150 ns,
'1' after 292950 ns, '0' after 293000 ns,
'1' after 303800 ns, '0' after 303850 ns,
'1' after 314650 ns, '0' after 314700 ns,
'1' after 325500 ns, '0' after 325550 ns,
'1' after 336350 ns, '0' after 336400 ns,
'1' after 347200 ns, '0' after 347250 ns,
'1' after 358050 ns, '0' after 358100 ns,
'1' after 368900 ns, '0' after 368950 ns,
'1' after 379750 ns, '0' after 379800 ns,
'1' after 390600 ns, '0' after 390650 ns,
'1' after 401450 ns, '0' after 401500 ns,
'1' after 412300 ns, '0' after 412350 ns,
'1' after 423150 ns, '0' after 423200 ns,
'1' after 434000 ns, '0' after 434050 ns,
'1' after 444850 ns, '0' after 444900 ns,
'1' after 455700 ns, '0' after 455750 ns,
'1' after 466550 ns, '0' after 466600 ns,
'1' after 477400 ns, '0' after 477450 ns,
'1' after 488250 ns, '0' after 488300 ns,
'1' after 499100 ns, '0' after 499150 ns,
'1' after 509950 ns, '0' after 510000 ns,
'1' after 520800 ns, '0' after 520850 ns,
'1' after 531650 ns, '0' after 531700 ns,
'1' after 542500 ns, '0' after 542550 ns,
'1' after 553350 ns, '0' after 553400 ns,
'1' after 564200 ns, '0' after 564250 ns,
'1' after 575050 ns, '0' after 575100 ns,
'1' after 585900 ns, '0' after 585950 ns,
'1' after 596750 ns, '0' after 596800 ns,
'1' after 607600 ns, '0' after 607650 ns,
'1' after 618450 ns, '0' after 618500 ns,
'1' after 629300 ns, '0' after 629350 ns,
'1' after 640150 ns, '0' after 640200 ns,
'1' after 651000 ns, '0' after 651050 ns,
'1' after 661850 ns, '0' after 661900 ns,
'1' after 672700 ns, '0' after 672750 ns,
'1' after 683550 ns, '0' after 683600 ns,
'1' after 694400 ns, '0' after 694450 ns,
'1' after 705250 ns, '0' after 705300 ns,
'1' after 716100 ns, '0' after 716150 ns,
'1' after 726950 ns, '0' after 727000 ns,
'1' after 737800 ns, '0' after 737850 ns,
'1' after 748650 ns, '0' after 748700 ns,
'1' after 759500 ns, '0' after 759550 ns,
'1' after 770350 ns, '0' after 770400 ns,
'1' after 781200 ns, '0' after 781250 ns,
'1' after 792050 ns, '0' after 792100 ns,
'1' after 802900 ns, '0' after 802950 ns,
'1' after 813750 ns, '0' after 813800 ns,
'1' after 824600 ns, '0' after 824650 ns,
'1' after 835450 ns, '0' after 835500 ns,
'1' after 846300 ns, '0' after 846350 ns,
'1' after 857150 ns, '0' after 857200 ns,
'1' after 868000 ns, '0' after 868050 ns,
'1' after 878850 ns, '0' after 878900 ns,
'1' after 889700 ns, '0' after 889750 ns,
'1' after 900550 ns, '0' after 900600 ns,
'1' after 911400 ns, '0' after 911450 ns,
'1' after 922250 ns, '0' after 922300 ns,
'1' after 933100 ns, '0' after 933150 ns,
'1' after 943950 ns, '0' after 944000 ns,
'1' after 954800 ns, '0' after 954850 ns,
'1' after 965650 ns, '0' after 965700 ns,
'1' after 976500 ns, '0' after 976550 ns,
'1' after 987350 ns, '0' after 987400 ns,
'1' after 998200 ns, '0' after 998250 ns,
'1' after 1009050 ns, '0' after 1009100 ns,
'1' after 1019900 ns, '0' after 1019950 ns,
'1' after 1030750 ns, '0' after 1030800 ns,
'1' after 1041600 ns, '0' after 1041650 ns,
'1' after 1052450 ns, '0' after 1052500 ns,
'1' after 1063300 ns, '0' after 1063350 ns,
'1' after 1074150 ns, '0' after 1074200 ns,
'1' after 1085000 ns, '0' after 1085050 ns,
'1' after 1095850 ns, '0' after 1095900 ns,
'1' after 1106700 ns, '0' after 1106750 ns,
'1' after 1117550 ns, '0' after 1117600 ns,
'1' after 1128400 ns, '0' after 1128450 ns,
'1' after 1139250 ns, '0' after 1139300 ns,
'1' after 1150100 ns, '0' after 1150150 ns,
'1' after 1160950 ns, '0' after 1161000 ns,
'1' after 1171800 ns, '0' after 1171850 ns,
'1' after 1182650 ns, '0' after 1182700 ns,
'1' after 1193500 ns, '0' after 1193550 ns,
'1' after 1204350 ns, '0' after 1204400 ns,
'1' after 1215200 ns, '0' after 1215250 ns,
'1' after 1226050 ns, '0' after 1226100 ns,
'1' after 1236900 ns, '0' after 1236950 ns,
'1' after 1247750 ns, '0' after 1247800 ns,
'1' after 1258600 ns, '0' after 1258650 ns,
'1' after 1269450 ns, '0' after 1269500 ns,
'1' after 1280300 ns, '0' after 1280350 ns,
'1' after 1291150 ns, '0' after 1291200 ns,
'1' after 1302000 ns, '0' after 1302050 ns,
'1' after 1312850 ns, '0' after 1312900 ns,
'1' after 1323700 ns, '0' after 1323750 ns,
'1' after 1334550 ns, '0' after 1334600 ns,
'1' after 1345400 ns, '0' after 1345450 ns,
'1' after 1356250 ns, '0' after 1356300 ns,
'1' after 1367100 ns, '0' after 1367150 ns,
'1' after 1377950 ns, '0' after 1378000 ns,
'1' after 1388800 ns, '0' after 1388850 ns,
'1' after 1399650 ns, '0' after 1399700 ns,
'1' after 1410500 ns, '0' after 1410550 ns,
'1' after 1421350 ns, '0' after 1421400 ns,
'1' after 1432200 ns, '0' after 1432250 ns,
'1' after 1443050 ns, '0' after 1443100 ns,
'1' after 1453900 ns, '0' after 1453950 ns,
'1' after 1464750 ns, '0' after 1464800 ns,
'1' after 1475600 ns, '0' after 1475650 ns,
'1' after 1486450 ns, '0' after 1486500 ns,
'1' after 1497300 ns, '0' after 1497350 ns,
'1' after 1508150 ns, '0' after 1508200 ns,
'1' after 1519000 ns, '0' after 1519050 ns,
'1' after 1529850 ns, '0' after 1529900 ns,
'1' after 1540700 ns, '0' after 1540750 ns,
'1' after 1551550 ns, '0' after 1551600 ns,
'1' after 1562400 ns, '0' after 1562450 ns,
'1' after 1573250 ns, '0' after 1573300 ns,
'1' after 1584100 ns, '0' after 1584150 ns,
'1' after 1594950 ns, '0' after 1595000 ns,
'1' after 1605800 ns, '0' after 1605850 ns,
'1' after 1616650 ns, '0' after 1616700 ns,
'1' after 1627500 ns, '0' after 1627550 ns,
'1' after 1638350 ns, '0' after 1638400 ns,
'1' after 1649200 ns, '0' after 1649250 ns,
'1' after 1660050 ns, '0' after 1660100 ns,
'1' after 1670900 ns, '0' after 1670950 ns,
'1' after 1681750 ns, '0' after 1681800 ns,
'1' after 1692600 ns, '0' after 1692650 ns,
'1' after 1703450 ns, '0' after 1703500 ns,
'1' after 1714300 ns, '0' after 1714350 ns,
'1' after 1725150 ns, '0' after 1725200 ns,
'1' after 1736000 ns, '0' after 1736050 ns,
'1' after 1746850 ns, '0' after 1746900 ns,
'1' after 1757700 ns, '0' after 1757750 ns,
'1' after 1768550 ns, '0' after 1768600 ns,
'1' after 1779400 ns, '0' after 1779450 ns,
'1' after 1790250 ns, '0' after 1790300 ns,
'1' after 1801100 ns, '0' after 1801150 ns,
'1' after 1811950 ns, '0' after 1812000 ns,
'1' after 1822800 ns, '0' after 1822850 ns,
'1' after 1833650 ns, '0' after 1833700 ns,
'1' after 1844500 ns, '0' after 1844550 ns,
'1' after 1855350 ns, '0' after 1855400 ns,
'1' after 1866200 ns, '0' after 1866250 ns,
'1' after 1877050 ns, '0' after 1877100 ns,
'1' after 1887900 ns, '0' after 1887950 ns,
'1' after 1898750 ns, '0' after 1898800 ns,
'1' after 1909600 ns, '0' after 1909650 ns,
'1' after 1920450 ns, '0' after 1920500 ns,
'1' after 1931300 ns, '0' after 1931350 ns,
'1' after 1942150 ns, '0' after 1942200 ns,
'1' after 1953000 ns, '0' after 1953050 ns,
'1' after 1963850 ns, '0' after 1963900 ns,
'1' after 1974700 ns, '0' after 1974750 ns,
'1' after 1985550 ns, '0' after 1985600 ns,
'1' after 1996400 ns, '0' after 1996450 ns,
'1' after 2007250 ns, '0' after 2007300 ns,
'1' after 2018100 ns, '0' after 2018150 ns,
'1' after 2028950 ns, '0' after 2029000 ns,
'1' after 2039800 ns, '0' after 2039850 ns,
'1' after 2050650 ns, '0' after 2050700 ns,
'1' after 2061500 ns, '0' after 2061550 ns,
'1' after 2072350 ns, '0' after 2072400 ns,
'1' after 2083200 ns, '0' after 2083250 ns,
'1' after 2094050 ns, '0' after 2094100 ns,
'1' after 2104900 ns, '0' after 2104950 ns,
'1' after 2115750 ns, '0' after 2115800 ns,
'1' after 2126600 ns, '0' after 2126650 ns,
'1' after 2137450 ns, '0' after 2137500 ns,
'1' after 2148300 ns, '0' after 2148350 ns,
'1' after 2159150 ns, '0' after 2159200 ns,
'1' after 2170000 ns, '0' after 2170050 ns,
'1' after 2180850 ns, '0' after 2180900 ns,
'1' after 2191700 ns, '0' after 2191750 ns,
'1' after 2202550 ns, '0' after 2202600 ns,
'1' after 2213400 ns, '0' after 2213450 ns,
'1' after 2224250 ns, '0' after 2224300 ns,
'1' after 2235100 ns, '0' after 2235150 ns,
'1' after 2245950 ns, '0' after 2246000 ns,
'1' after 2256800 ns, '0' after 2256850 ns,
'1' after 2267650 ns, '0' after 2267700 ns,
'1' after 2278500 ns, '0' after 2278550 ns,
'1' after 2289350 ns, '0' after 2289400 ns,
'1' after 2300200 ns, '0' after 2300250 ns,
'1' after 2311050 ns, '0' after 2311100 ns,
'1' after 2321900 ns, '0' after 2321950 ns,
'1' after 2332750 ns, '0' after 2332800 ns,
'1' after 2343600 ns, '0' after 2343650 ns,
'1' after 2354450 ns, '0' after 2354500 ns,
'1' after 2365300 ns, '0' after 2365350 ns,
'1' after 2376150 ns, '0' after 2376200 ns,
'1' after 2387000 ns, '0' after 2387050 ns,
'1' after 2397850 ns, '0' after 2397900 ns,
'1' after 2408700 ns, '0' after 2408750 ns,
'1' after 2419550 ns, '0' after 2419600 ns,
'1' after 2430400 ns, '0' after 2430450 ns,
'1' after 2441250 ns, '0' after 2441300 ns,
'1' after 2452100 ns, '0' after 2452150 ns,
'1' after 2462950 ns, '0' after 2463000 ns,
'1' after 2473800 ns, '0' after 2473850 ns,
'1' after 2484650 ns, '0' after 2484700 ns,
'1' after 2495500 ns, '0' after 2495550 ns,
'1' after 2506350 ns, '0' after 2506400 ns,
'1' after 2517200 ns, '0' after 2517250 ns,
'1' after 2528050 ns, '0' after 2528100 ns,
'1' after 2538900 ns, '0' after 2538950 ns,
'1' after 2549750 ns, '0' after 2549800 ns,
'1' after 2560600 ns, '0' after 2560650 ns,
'1' after 2571450 ns, '0' after 2571500 ns,
'1' after 2582300 ns, '0' after 2582350 ns,
'1' after 2593150 ns, '0' after 2593200 ns,
'1' after 2604000 ns, '0' after 2604050 ns,
'1' after 2614850 ns, '0' after 2614900 ns,
'1' after 2625700 ns, '0' after 2625750 ns,
'1' after 2636550 ns, '0' after 2636600 ns,
'1' after 2647400 ns, '0' after 2647450 ns,
'1' after 2658250 ns, '0' after 2658300 ns,
'1' after 2669100 ns, '0' after 2669150 ns,
'1' after 2679950 ns, '0' after 2680000 ns,
'1' after 2690800 ns, '0' after 2690850 ns,
'1' after 2701650 ns, '0' after 2701700 ns,
'1' after 2712500 ns, '0' after 2712550 ns,
'1' after 2723350 ns, '0' after 2723400 ns,
'1' after 2734200 ns, '0' after 2734250 ns,
'1' after 2745050 ns, '0' after 2745100 ns,
'1' after 2755900 ns, '0' after 2755950 ns,
'1' after 2766750 ns, '0' after 2766800 ns,
'1' after 2777600 ns, '0' after 2777650 ns,
'1' after 2788450 ns, '0' after 2788500 ns,
'1' after 2799300 ns, '0' after 2799350 ns,
'1' after 2810150 ns, '0' after 2810200 ns,
'1' after 2821000 ns, '0' after 2821050 ns,
'1' after 2831850 ns, '0' after 2831900 ns,
'1' after 2842700 ns, '0' after 2842750 ns,
'1' after 2853550 ns, '0' after 2853600 ns,
'1' after 2864400 ns, '0' after 2864450 ns,
'1' after 2875250 ns, '0' after 2875300 ns,
'1' after 2886100 ns, '0' after 2886150 ns,
'1' after 2896950 ns, '0' after 2897000 ns,
'1' after 2907800 ns, '0' after 2907850 ns,
'1' after 2918650 ns, '0' after 2918700 ns,
'1' after 2929500 ns, '0' after 2929550 ns,
'1' after 2940350 ns, '0' after 2940400 ns,
'1' after 2951200 ns, '0' after 2951250 ns,
'1' after 2962050 ns, '0' after 2962100 ns,
'1' after 2972900 ns, '0' after 2972950 ns,
'1' after 2983750 ns, '0' after 2983800 ns,
'1' after 2994600 ns, '0' after 2994650 ns,
'1' after 3005450 ns, '0' after 3005500 ns,
'1' after 3016300 ns, '0' after 3016350 ns,
'1' after 3027150 ns, '0' after 3027200 ns,
'1' after 3038000 ns, '0' after 3038050 ns,
'1' after 3048850 ns, '0' after 3048900 ns,
'1' after 3059700 ns, '0' after 3059750 ns,
'1' after 3070550 ns, '0' after 3070600 ns,
'1' after 3081400 ns, '0' after 3081450 ns,
'1' after 3092250 ns, '0' after 3092300 ns,
'1' after 3103100 ns, '0' after 3103150 ns,
'1' after 3113950 ns, '0' after 3114000 ns,
'1' after 3124800 ns, '0' after 3124850 ns,
'1' after 3135650 ns, '0' after 3135700 ns,
'1' after 3146500 ns, '0' after 3146550 ns,
'1' after 3157350 ns, '0' after 3157400 ns,
'1' after 3168200 ns, '0' after 3168250 ns,
'1' after 3179050 ns, '0' after 3179100 ns,
'1' after 3189900 ns, '0' after 3189950 ns,
'1' after 3200750 ns, '0' after 3200800 ns,
'1' after 3211600 ns, '0' after 3211650 ns,
'1' after 3222450 ns, '0' after 3222500 ns,
'1' after 3233300 ns, '0' after 3233350 ns,
'1' after 3244150 ns, '0' after 3244200 ns,
'1' after 3255000 ns, '0' after 3255050 ns,
'1' after 3265850 ns, '0' after 3265900 ns,
'1' after 3276700 ns, '0' after 3276750 ns,
'1' after 3287550 ns, '0' after 3287600 ns,
'1' after 3298400 ns, '0' after 3298450 ns,
'1' after 3309250 ns, '0' after 3309300 ns,
'1' after 3320100 ns, '0' after 3320150 ns,
'1' after 3330950 ns, '0' after 3331000 ns,
'1' after 3341800 ns, '0' after 3341850 ns,
'1' after 3352650 ns, '0' after 3352700 ns,
'1' after 3363500 ns, '0' after 3363550 ns,
'1' after 3374350 ns, '0' after 3374400 ns,
'1' after 3385200 ns, '0' after 3385250 ns,
'1' after 3396050 ns, '0' after 3396100 ns,
'1' after 3406900 ns, '0' after 3406950 ns,
'1' after 3417750 ns, '0' after 3417800 ns,
'1' after 3428600 ns, '0' after 3428650 ns,
'1' after 3439450 ns, '0' after 3439500 ns,
'1' after 3450300 ns, '0' after 3450350 ns,
'1' after 3461150 ns, '0' after 3461200 ns,
'1' after 3472000 ns, '0' after 3472050 ns,
'1' after 3482850 ns, '0' after 3482900 ns,
'1' after 3493700 ns, '0' after 3493750 ns,
'1' after 3504550 ns, '0' after 3504600 ns,
'1' after 3515400 ns, '0' after 3515450 ns,
'1' after 3526250 ns, '0' after 3526300 ns,
'1' after 3537100 ns, '0' after 3537150 ns,
'1' after 3547950 ns, '0' after 3548000 ns,
'1' after 3558800 ns, '0' after 3558850 ns,
'1' after 3569650 ns, '0' after 3569700 ns,
'1' after 3580500 ns, '0' after 3580550 ns,
'1' after 3591350 ns, '0' after 3591400 ns,
'1' after 3602200 ns, '0' after 3602250 ns,
'1' after 3613050 ns, '0' after 3613100 ns,
'1' after 3623900 ns, '0' after 3623950 ns,
'1' after 3634750 ns, '0' after 3634800 ns,
'1' after 3645600 ns, '0' after 3645650 ns,
'1' after 3656450 ns, '0' after 3656500 ns,
'1' after 3667300 ns, '0' after 3667350 ns,
'1' after 3678150 ns, '0' after 3678200 ns,
'1' after 3689000 ns, '0' after 3689050 ns,
'1' after 3699850 ns, '0' after 3699900 ns,
'1' after 3710700 ns, '0' after 3710750 ns,
'1' after 3721550 ns, '0' after 3721600 ns,
'1' after 3732400 ns, '0' after 3732450 ns,
'1' after 3743250 ns, '0' after 3743300 ns,
'1' after 3754100 ns, '0' after 3754150 ns,
'1' after 3764950 ns, '0' after 3765000 ns,
'1' after 3775800 ns, '0' after 3775850 ns,
'1' after 3786650 ns, '0' after 3786700 ns,
'1' after 3797500 ns, '0' after 3797550 ns,
'1' after 3808350 ns, '0' after 3808400 ns,
'1' after 3819200 ns, '0' after 3819250 ns,
'1' after 3830050 ns, '0' after 3830100 ns,
'1' after 3840900 ns, '0' after 3840950 ns,
'1' after 3851750 ns, '0' after 3851800 ns,
'1' after 3862600 ns, '0' after 3862650 ns,
'1' after 3873450 ns, '0' after 3873500 ns,
'1' after 3884300 ns, '0' after 3884350 ns,
'1' after 3895150 ns, '0' after 3895200 ns,
'1' after 3906000 ns, '0' after 3906050 ns,
'1' after 3916850 ns, '0' after 3916900 ns,
'1' after 3927700 ns, '0' after 3927750 ns,
'1' after 3938550 ns, '0' after 3938600 ns,
'1' after 3949400 ns, '0' after 3949450 ns,
'1' after 3960250 ns, '0' after 3960300 ns,
'1' after 3971100 ns, '0' after 3971150 ns,
'1' after 3981950 ns, '0' after 3982000 ns,
'1' after 3992800 ns, '0' after 3992850 ns,
'1' after 4003650 ns, '0' after 4003700 ns,
'1' after 4014500 ns, '0' after 4014550 ns,
'1' after 4025350 ns, '0' after 4025400 ns,
'1' after 4036200 ns, '0' after 4036250 ns,
'1' after 4047050 ns, '0' after 4047100 ns,
'1' after 4057900 ns, '0' after 4057950 ns,
'1' after 4068750 ns, '0' after 4068800 ns,
'1' after 4079600 ns, '0' after 4079650 ns,
'1' after 4090450 ns, '0' after 4090500 ns,
'1' after 4101300 ns, '0' after 4101350 ns,
'1' after 4112150 ns, '0' after 4112200 ns,
'1' after 4123000 ns, '0' after 4123050 ns,
'1' after 4133850 ns, '0' after 4133900 ns,
'1' after 4144700 ns, '0' after 4144750 ns,
'1' after 4155550 ns, '0' after 4155600 ns,
'1' after 4166400 ns, '0' after 4166450 ns,
'1' after 4177250 ns, '0' after 4177300 ns,
'1' after 4188100 ns, '0' after 4188150 ns,
'1' after 4198950 ns, '0' after 4199000 ns,
'1' after 4209800 ns, '0' after 4209850 ns,
'1' after 4220650 ns, '0' after 4220700 ns,
'1' after 4231500 ns, '0' after 4231550 ns,
'1' after 4242350 ns, '0' after 4242400 ns,
'1' after 4253200 ns, '0' after 4253250 ns,
'1' after 4264050 ns, '0' after 4264100 ns,
'1' after 4274900 ns, '0' after 4274950 ns,
'1' after 4285750 ns, '0' after 4285800 ns,
'1' after 4296600 ns, '0' after 4296650 ns,
'1' after 4307450 ns, '0' after 4307500 ns,
'1' after 4318300 ns, '0' after 4318350 ns,
'1' after 4329150 ns, '0' after 4329200 ns,
'1' after 4340000 ns, '0' after 4340050 ns,
'1' after 4350850 ns, '0' after 4350900 ns,
'1' after 4361700 ns, '0' after 4361750 ns,
'1' after 4372550 ns, '0' after 4372600 ns,
'1' after 4383400 ns, '0' after 4383450 ns,
'1' after 4394250 ns, '0' after 4394300 ns,
'1' after 4405100 ns, '0' after 4405150 ns,
'1' after 4415950 ns, '0' after 4416000 ns,
'1' after 4426800 ns, '0' after 4426850 ns,
'1' after 4437650 ns, '0' after 4437700 ns,
'1' after 4448500 ns, '0' after 4448550 ns,
'1' after 4459350 ns, '0' after 4459400 ns,
'1' after 4470200 ns, '0' after 4470250 ns,
'1' after 4481050 ns, '0' after 4481100 ns,
'1' after 4491900 ns, '0' after 4491950 ns,
'1' after 4502750 ns, '0' after 4502800 ns,
'1' after 4513600 ns, '0' after 4513650 ns,
'1' after 4524450 ns, '0' after 4524500 ns,
'1' after 4535300 ns, '0' after 4535350 ns,
'1' after 4546150 ns, '0' after 4546200 ns,
'1' after 4557000 ns, '0' after 4557050 ns,
'1' after 4567850 ns, '0' after 4567900 ns,
'1' after 4578700 ns, '0' after 4578750 ns,
'1' after 4589550 ns, '0' after 4589600 ns,
'1' after 4600400 ns, '0' after 4600450 ns,
'1' after 4611250 ns, '0' after 4611300 ns,
'1' after 4622100 ns, '0' after 4622150 ns,
'1' after 4632950 ns, '0' after 4633000 ns,
'1' after 4643800 ns, '0' after 4643850 ns,
'1' after 4654650 ns, '0' after 4654700 ns,
'1' after 4665500 ns, '0' after 4665550 ns,
'1' after 4676350 ns, '0' after 4676400 ns,
'1' after 4687200 ns, '0' after 4687250 ns,
'1' after 4698050 ns, '0' after 4698100 ns,
'1' after 4708900 ns, '0' after 4708950 ns,
'1' after 4719750 ns, '0' after 4719800 ns,
'1' after 4730600 ns, '0' after 4730650 ns,
'1' after 4741450 ns, '0' after 4741500 ns,
'1' after 4752300 ns, '0' after 4752350 ns,
'1' after 4763150 ns, '0' after 4763200 ns,
'1' after 4774000 ns, '0' after 4774050 ns,
'1' after 4784850 ns, '0' after 4784900 ns,
'1' after 4795700 ns, '0' after 4795750 ns,
'1' after 4806550 ns, '0' after 4806600 ns,
'1' after 4817400 ns, '0' after 4817450 ns,
'1' after 4828250 ns, '0' after 4828300 ns,
'1' after 4839100 ns, '0' after 4839150 ns,
'1' after 4849950 ns, '0' after 4850000 ns,
'1' after 4860800 ns, '0' after 4860850 ns,
'1' after 4871650 ns, '0' after 4871700 ns,
'1' after 4882500 ns, '0' after 4882550 ns,
'1' after 4893350 ns, '0' after 4893400 ns,
'1' after 4904200 ns, '0' after 4904250 ns,
'1' after 4915050 ns, '0' after 4915100 ns,
'1' after 4925900 ns, '0' after 4925950 ns,
'1' after 4936750 ns, '0' after 4936800 ns,
'1' after 4947600 ns, '0' after 4947650 ns,
'1' after 4958450 ns, '0' after 4958500 ns,
'1' after 4969300 ns, '0' after 4969350 ns,
'1' after 4980150 ns, '0' after 4980200 ns,
'1' after 4991000 ns, '0' after 4991050 ns,
'1' after 5001850 ns, '0' after 5001900 ns,
'1' after 5012700 ns, '0' after 5012750 ns,
'1' after 5023550 ns, '0' after 5023600 ns,
'1' after 5034400 ns, '0' after 5034450 ns,
'1' after 5045250 ns, '0' after 5045300 ns,
'1' after 5056100 ns, '0' after 5056150 ns,
'1' after 5066950 ns, '0' after 5067000 ns,
'1' after 5077800 ns, '0' after 5077850 ns,
'1' after 5088650 ns, '0' after 5088700 ns,
'1' after 5099500 ns, '0' after 5099550 ns,
'1' after 5110350 ns, '0' after 5110400 ns,
'1' after 5121200 ns, '0' after 5121250 ns,
'1' after 5132050 ns, '0' after 5132100 ns,
'1' after 5142900 ns, '0' after 5142950 ns,
'1' after 5153750 ns, '0' after 5153800 ns,
'1' after 5164600 ns, '0' after 5164650 ns,
'1' after 5175450 ns, '0' after 5175500 ns,
'1' after 5186300 ns, '0' after 5186350 ns,
'1' after 5197150 ns, '0' after 5197200 ns,
'1' after 5208000 ns, '0' after 5208050 ns,
'1' after 5218850 ns, '0' after 5218900 ns,
'1' after 5229700 ns, '0' after 5229750 ns,
'1' after 5240550 ns, '0' after 5240600 ns,
'1' after 5251400 ns, '0' after 5251450 ns,
'1' after 5262250 ns, '0' after 5262300 ns,
'1' after 5273100 ns, '0' after 5273150 ns,
'1' after 5283950 ns, '0' after 5284000 ns,
'1' after 5294800 ns, '0' after 5294850 ns,
'1' after 5305650 ns, '0' after 5305700 ns,
'1' after 5316500 ns, '0' after 5316550 ns,
'1' after 5327350 ns, '0' after 5327400 ns,
'1' after 5338200 ns, '0' after 5338250 ns,
'1' after 5349050 ns, '0' after 5349100 ns,
'1' after 5359900 ns, '0' after 5359950 ns,
'1' after 5370750 ns, '0' after 5370800 ns,
'1' after 5381600 ns, '0' after 5381650 ns,
'1' after 5392450 ns, '0' after 5392500 ns,
'1' after 5403300 ns, '0' after 5403350 ns,
'1' after 5414150 ns, '0' after 5414200 ns,
'1' after 5425000 ns, '0' after 5425050 ns,
'1' after 5435850 ns, '0' after 5435900 ns,
'1' after 5446700 ns, '0' after 5446750 ns,
'1' after 5457550 ns, '0' after 5457600 ns,
'1' after 5468400 ns, '0' after 5468450 ns,
'1' after 5479250 ns, '0' after 5479300 ns,
'1' after 5490100 ns, '0' after 5490150 ns,
'1' after 5500950 ns, '0' after 5501000 ns,
'1' after 5511800 ns, '0' after 5511850 ns,
'1' after 5522650 ns, '0' after 5522700 ns,
'1' after 5533500 ns, '0' after 5533550 ns,
'1' after 5544350 ns, '0' after 5544400 ns,
'1' after 5555200 ns, '0' after 5555250 ns,
'1' after 5566050 ns, '0' after 5566100 ns,
'1' after 5576900 ns, '0' after 5576950 ns,
'1' after 5587750 ns, '0' after 5587800 ns,
'1' after 5598600 ns, '0' after 5598650 ns,
'1' after 5609450 ns, '0' after 5609500 ns,
'1' after 5620300 ns, '0' after 5620350 ns,
'1' after 5631150 ns, '0' after 5631200 ns,
'1' after 5642000 ns, '0' after 5642050 ns,
'1' after 5652850 ns, '0' after 5652900 ns,
'1' after 5663700 ns, '0' after 5663750 ns,
'1' after 5674550 ns, '0' after 5674600 ns,
'1' after 5685400 ns, '0' after 5685450 ns,
'1' after 5696250 ns, '0' after 5696300 ns,
'1' after 5707100 ns, '0' after 5707150 ns,
'1' after 5717950 ns, '0' after 5718000 ns,
'1' after 5728800 ns, '0' after 5728850 ns,
'1' after 5739650 ns, '0' after 5739700 ns,
'1' after 5750500 ns, '0' after 5750550 ns,
'1' after 5761350 ns, '0' after 5761400 ns,
'1' after 5772200 ns, '0' after 5772250 ns,
'1' after 5783050 ns, '0' after 5783100 ns,
'1' after 5793900 ns, '0' after 5793950 ns,
'1' after 5804750 ns, '0' after 5804800 ns,
'1' after 5815600 ns, '0' after 5815650 ns,
'1' after 5826450 ns, '0' after 5826500 ns,
'1' after 5837300 ns, '0' after 5837350 ns,
'1' after 5848150 ns, '0' after 5848200 ns,
'1' after 5859000 ns, '0' after 5859050 ns,
'1' after 5869850 ns, '0' after 5869900 ns,
'1' after 5880700 ns, '0' after 5880750 ns,
'1' after 5891550 ns, '0' after 5891600 ns,
'1' after 5902400 ns, '0' after 5902450 ns,
'1' after 5913250 ns, '0' after 5913300 ns,
'1' after 5924100 ns, '0' after 5924150 ns,
'1' after 5934950 ns, '0' after 5935000 ns,
'1' after 5945800 ns, '0' after 5945850 ns,
'1' after 5956650 ns, '0' after 5956700 ns,
'1' after 5967500 ns, '0' after 5967550 ns,
'1' after 5978350 ns, '0' after 5978400 ns,
'1' after 5989200 ns, '0' after 5989250 ns,
'1' after 6000050 ns, '0' after 6000100 ns,
'1' after 6010900 ns, '0' after 6010950 ns,
'1' after 6021750 ns, '0' after 6021800 ns,
'1' after 6032600 ns, '0' after 6032650 ns,
'1' after 6043450 ns, '0' after 6043500 ns,
'1' after 6054300 ns, '0' after 6054350 ns,
'1' after 6065150 ns, '0' after 6065200 ns,
'1' after 6076000 ns, '0' after 6076050 ns,
'1' after 6086850 ns, '0' after 6086900 ns,
'1' after 6097700 ns, '0' after 6097750 ns,
'1' after 6108550 ns, '0' after 6108600 ns,
'1' after 6119400 ns, '0' after 6119450 ns,
'1' after 6130250 ns, '0' after 6130300 ns,
'1' after 6141100 ns, '0' after 6141150 ns,
'1' after 6151950 ns, '0' after 6152000 ns,
'1' after 6162800 ns, '0' after 6162850 ns,
'1' after 6173650 ns, '0' after 6173700 ns,
'1' after 6184500 ns, '0' after 6184550 ns,
'1' after 6195350 ns, '0' after 6195400 ns,
'1' after 6206200 ns, '0' after 6206250 ns,
'1' after 6217050 ns, '0' after 6217100 ns,
'1' after 6227900 ns, '0' after 6227950 ns,
'1' after 6238750 ns, '0' after 6238800 ns,
'1' after 6249600 ns, '0' after 6249650 ns,
'1' after 6260450 ns, '0' after 6260500 ns,
'1' after 6271300 ns, '0' after 6271350 ns,
'1' after 6282150 ns, '0' after 6282200 ns,
'1' after 6293000 ns, '0' after 6293050 ns,
'1' after 6303850 ns, '0' after 6303900 ns,
'1' after 6314700 ns, '0' after 6314750 ns,
'1' after 6325550 ns, '0' after 6325600 ns,
'1' after 6336400 ns, '0' after 6336450 ns,
'1' after 6347250 ns, '0' after 6347300 ns,
'1' after 6358100 ns, '0' after 6358150 ns,
'1' after 6368950 ns, '0' after 6369000 ns,
'1' after 6379800 ns, '0' after 6379850 ns,
'1' after 6390650 ns, '0' after 6390700 ns,
'1' after 6401500 ns, '0' after 6401550 ns,
'1' after 6412350 ns, '0' after 6412400 ns,
'1' after 6423200 ns, '0' after 6423250 ns,
'1' after 6434050 ns, '0' after 6434100 ns,
'1' after 6444900 ns, '0' after 6444950 ns,
'1' after 6455750 ns, '0' after 6455800 ns,
'1' after 6466600 ns, '0' after 6466650 ns,
'1' after 6477450 ns, '0' after 6477500 ns,
'1' after 6488300 ns, '0' after 6488350 ns,
'1' after 6499150 ns, '0' after 6499200 ns,
'1' after 6510000 ns, '0' after 6510050 ns,
'1' after 6520850 ns, '0' after 6520900 ns,
'1' after 6531700 ns, '0' after 6531750 ns,
'1' after 6542550 ns, '0' after 6542600 ns,
'1' after 6553400 ns, '0' after 6553450 ns,
'1' after 6564250 ns, '0' after 6564300 ns,
'1' after 6575100 ns, '0' after 6575150 ns,
'1' after 6585950 ns, '0' after 6586000 ns,
'1' after 6596800 ns, '0' after 6596850 ns,
'1' after 6607650 ns, '0' after 6607700 ns,
'1' after 6618500 ns, '0' after 6618550 ns,
'1' after 6629350 ns, '0' after 6629400 ns,
'1' after 6640200 ns, '0' after 6640250 ns,
'1' after 6651050 ns, '0' after 6651100 ns,
'1' after 6661900 ns, '0' after 6661950 ns,
'1' after 6672750 ns, '0' after 6672800 ns,
'1' after 6683600 ns, '0' after 6683650 ns,
'1' after 6694450 ns, '0' after 6694500 ns,
'1' after 6705300 ns, '0' after 6705350 ns,
'1' after 6716150 ns, '0' after 6716200 ns,
'1' after 6727000 ns, '0' after 6727050 ns,
'1' after 6737850 ns, '0' after 6737900 ns,
'1' after 6748700 ns, '0' after 6748750 ns,
'1' after 6759550 ns, '0' after 6759600 ns,
'1' after 6770400 ns, '0' after 6770450 ns,
'1' after 6781250 ns, '0' after 6781300 ns,
'1' after 6792100 ns, '0' after 6792150 ns,
'1' after 6802950 ns, '0' after 6803000 ns,
'1' after 6813800 ns, '0' after 6813850 ns,
'1' after 6824650 ns, '0' after 6824700 ns,
'1' after 6835500 ns, '0' after 6835550 ns,
'1' after 6846350 ns, '0' after 6846400 ns,
'1' after 6857200 ns, '0' after 6857250 ns,
'1' after 6868050 ns, '0' after 6868100 ns,
'1' after 6878900 ns, '0' after 6878950 ns,
'1' after 6889750 ns, '0' after 6889800 ns,
'1' after 6900600 ns, '0' after 6900650 ns,
'1' after 6911450 ns, '0' after 6911500 ns,
'1' after 6922300 ns, '0' after 6922350 ns,
'1' after 6933150 ns, '0' after 6933200 ns,
'1' after 6944000 ns, '0' after 6944050 ns,
'1' after 6954850 ns, '0' after 6954900 ns,
'1' after 6965700 ns, '0' after 6965750 ns,
'1' after 6976550 ns, '0' after 6976600 ns,
'1' after 6987400 ns, '0' after 6987450 ns,
'1' after 6998250 ns, '0' after 6998300 ns,
'1' after 7009100 ns, '0' after 7009150 ns,
'1' after 7019950 ns, '0' after 7020000 ns,
'1' after 7030800 ns, '0' after 7030850 ns,
'1' after 7041650 ns, '0' after 7041700 ns,
'1' after 7052500 ns, '0' after 7052550 ns,
'1' after 7063350 ns, '0' after 7063400 ns,
'1' after 7074200 ns, '0' after 7074250 ns,
'1' after 7085050 ns, '0' after 7085100 ns,
'1' after 7095900 ns, '0' after 7095950 ns,
'1' after 7106750 ns, '0' after 7106800 ns,
'1' after 7117600 ns, '0' after 7117650 ns,
'1' after 7128450 ns, '0' after 7128500 ns,
'1' after 7139300 ns, '0' after 7139350 ns,
'1' after 7150150 ns, '0' after 7150200 ns,
'1' after 7161000 ns, '0' after 7161050 ns,
'1' after 7171850 ns, '0' after 7171900 ns,
'1' after 7182700 ns, '0' after 7182750 ns,
'1' after 7193550 ns, '0' after 7193600 ns,
'1' after 7204400 ns, '0' after 7204450 ns,
'1' after 7215250 ns, '0' after 7215300 ns,
'1' after 7226100 ns, '0' after 7226150 ns,
'1' after 7236950 ns, '0' after 7237000 ns,
'1' after 7247800 ns, '0' after 7247850 ns,
'1' after 7258650 ns, '0' after 7258700 ns,
'1' after 7269500 ns, '0' after 7269550 ns,
'1' after 7280350 ns, '0' after 7280400 ns,
'1' after 7291200 ns, '0' after 7291250 ns,
'1' after 7302050 ns, '0' after 7302100 ns,
'1' after 7312900 ns, '0' after 7312950 ns,
'1' after 7323750 ns, '0' after 7323800 ns,
'1' after 7334600 ns, '0' after 7334650 ns,
'1' after 7345450 ns, '0' after 7345500 ns,
'1' after 7356300 ns, '0' after 7356350 ns,
'1' after 7367150 ns, '0' after 7367200 ns,
'1' after 7378000 ns, '0' after 7378050 ns,
'1' after 7388850 ns, '0' after 7388900 ns,
'1' after 7399700 ns, '0' after 7399750 ns,
'1' after 7410550 ns, '0' after 7410600 ns,
'1' after 7421400 ns, '0' after 7421450 ns,
'1' after 7432250 ns, '0' after 7432300 ns,
'1' after 7443100 ns, '0' after 7443150 ns,
'1' after 7453950 ns, '0' after 7454000 ns,
'1' after 7464800 ns, '0' after 7464850 ns,
'1' after 7475650 ns, '0' after 7475700 ns,
'1' after 7486500 ns, '0' after 7486550 ns,
'1' after 7497350 ns, '0' after 7497400 ns,
'1' after 7508200 ns, '0' after 7508250 ns,
'1' after 7519050 ns, '0' after 7519100 ns,
'1' after 7529900 ns, '0' after 7529950 ns,
'1' after 7540750 ns, '0' after 7540800 ns,
'1' after 7551600 ns, '0' after 7551650 ns,
'1' after 7562450 ns, '0' after 7562500 ns,
'1' after 7573300 ns, '0' after 7573350 ns,
'1' after 7584150 ns, '0' after 7584200 ns,
'1' after 7595000 ns, '0' after 7595050 ns,
'1' after 7605850 ns, '0' after 7605900 ns,
'1' after 7616700 ns, '0' after 7616750 ns,
'1' after 7627550 ns, '0' after 7627600 ns,
'1' after 7638400 ns, '0' after 7638450 ns,
'1' after 7649250 ns, '0' after 7649300 ns,
'1' after 7660100 ns, '0' after 7660150 ns,
'1' after 7670950 ns, '0' after 7671000 ns,
'1' after 7681800 ns, '0' after 7681850 ns,
'1' after 7692650 ns, '0' after 7692700 ns,
'1' after 7703500 ns, '0' after 7703550 ns,
'1' after 7714350 ns, '0' after 7714400 ns,
'1' after 7725200 ns, '0' after 7725250 ns,
'1' after 7736050 ns, '0' after 7736100 ns,
'1' after 7746900 ns, '0' after 7746950 ns,
'1' after 7757750 ns, '0' after 7757800 ns,
'1' after 7768600 ns, '0' after 7768650 ns,
'1' after 7779450 ns, '0' after 7779500 ns,
'1' after 7790300 ns, '0' after 7790350 ns,
'1' after 7801150 ns, '0' after 7801200 ns,
'1' after 7812000 ns, '0' after 7812050 ns,
'1' after 7822850 ns, '0' after 7822900 ns,
'1' after 7833700 ns, '0' after 7833750 ns,
'1' after 7844550 ns, '0' after 7844600 ns,
'1' after 7855400 ns, '0' after 7855450 ns,
'1' after 7866250 ns, '0' after 7866300 ns,
'1' after 7877100 ns, '0' after 7877150 ns,
'1' after 7887950 ns, '0' after 7888000 ns,
'1' after 7898800 ns, '0' after 7898850 ns,
'1' after 7909650 ns, '0' after 7909700 ns,
'1' after 7920500 ns, '0' after 7920550 ns,
'1' after 7931350 ns, '0' after 7931400 ns,
'1' after 7942200 ns, '0' after 7942250 ns,
'1' after 7953050 ns, '0' after 7953100 ns,
'1' after 7963900 ns, '0' after 7963950 ns,
'1' after 7974750 ns, '0' after 7974800 ns,
'1' after 7985600 ns, '0' after 7985650 ns,
'1' after 7996450 ns, '0' after 7996500 ns,
'1' after 8007300 ns, '0' after 8007350 ns,
'1' after 8018150 ns, '0' after 8018200 ns,
'1' after 8029000 ns, '0' after 8029050 ns,
'1' after 8039850 ns, '0' after 8039900 ns,
'1' after 8050700 ns, '0' after 8050750 ns,
'1' after 8061550 ns, '0' after 8061600 ns,
'1' after 8072400 ns, '0' after 8072450 ns,
'1' after 8083250 ns, '0' after 8083300 ns,
'1' after 8094100 ns, '0' after 8094150 ns,
'1' after 8104950 ns, '0' after 8105000 ns,
'1' after 8115800 ns, '0' after 8115850 ns,
'1' after 8126650 ns, '0' after 8126700 ns,
'1' after 8137500 ns, '0' after 8137550 ns,
'1' after 8148350 ns, '0' after 8148400 ns,
'1' after 8159200 ns, '0' after 8159250 ns,
'1' after 8170050 ns, '0' after 8170100 ns,
'1' after 8180900 ns, '0' after 8180950 ns,
'1' after 8191750 ns, '0' after 8191800 ns,
'1' after 8202600 ns, '0' after 8202650 ns,
'1' after 8213450 ns, '0' after 8213500 ns,
'1' after 8224300 ns, '0' after 8224350 ns,
'1' after 8235150 ns, '0' after 8235200 ns,
'1' after 8246000 ns, '0' after 8246050 ns,
'1' after 8256850 ns, '0' after 8256900 ns,
'1' after 8267700 ns, '0' after 8267750 ns,
'1' after 8278550 ns, '0' after 8278600 ns,
'1' after 8289400 ns, '0' after 8289450 ns,
'1' after 8300250 ns, '0' after 8300300 ns,
'1' after 8311100 ns, '0' after 8311150 ns,
'1' after 8321950 ns, '0' after 8322000 ns,
'1' after 8332800 ns, '0' after 8332850 ns,
'1' after 8343650 ns, '0' after 8343700 ns,
'1' after 8354500 ns, '0' after 8354550 ns,
'1' after 8365350 ns, '0' after 8365400 ns,
'1' after 8376200 ns, '0' after 8376250 ns,
'1' after 8387050 ns, '0' after 8387100 ns,
'1' after 8397900 ns, '0' after 8397950 ns,
'1' after 8408750 ns, '0' after 8408800 ns,
'1' after 8419600 ns, '0' after 8419650 ns,
'1' after 8430450 ns, '0' after 8430500 ns,
'1' after 8441300 ns, '0' after 8441350 ns,
'1' after 8452150 ns, '0' after 8452200 ns,
'1' after 8463000 ns, '0' after 8463050 ns,
'1' after 8473850 ns, '0' after 8473900 ns,
'1' after 8484700 ns, '0' after 8484750 ns,
'1' after 8495550 ns, '0' after 8495600 ns,
'1' after 8506400 ns, '0' after 8506450 ns,
'1' after 8517250 ns, '0' after 8517300 ns,
'1' after 8528100 ns, '0' after 8528150 ns,
'1' after 8538950 ns, '0' after 8539000 ns,
'1' after 8549800 ns, '0' after 8549850 ns,
'1' after 8560650 ns, '0' after 8560700 ns,
'1' after 8571500 ns, '0' after 8571550 ns,
'1' after 8582350 ns, '0' after 8582400 ns,
'1' after 8593200 ns, '0' after 8593250 ns,
'1' after 8604050 ns, '0' after 8604100 ns,
'1' after 8614900 ns, '0' after 8614950 ns,
'1' after 8625750 ns, '0' after 8625800 ns,
'1' after 8636600 ns, '0' after 8636650 ns,
'1' after 8647450 ns, '0' after 8647500 ns,
'1' after 8658300 ns, '0' after 8658350 ns,
'1' after 8669150 ns, '0' after 8669200 ns,
'1' after 8680000 ns, '0' after 8680050 ns,
'1' after 8690850 ns, '0' after 8690900 ns,
'1' after 8701700 ns, '0' after 8701750 ns,
'1' after 8712550 ns, '0' after 8712600 ns,
'1' after 8723400 ns, '0' after 8723450 ns,
'1' after 8734250 ns, '0' after 8734300 ns,
'1' after 8745100 ns, '0' after 8745150 ns,
'1' after 8755950 ns, '0' after 8756000 ns,
'1' after 8766800 ns, '0' after 8766850 ns,
'1' after 8777650 ns, '0' after 8777700 ns,
'1' after 8788500 ns, '0' after 8788550 ns,
'1' after 8799350 ns, '0' after 8799400 ns,
'1' after 8810200 ns, '0' after 8810250 ns,
'1' after 8821050 ns, '0' after 8821100 ns,
'1' after 8831900 ns, '0' after 8831950 ns,
'1' after 8842750 ns, '0' after 8842800 ns,
'1' after 8853600 ns, '0' after 8853650 ns,
'1' after 8864450 ns, '0' after 8864500 ns,
'1' after 8875300 ns, '0' after 8875350 ns,
'1' after 8886150 ns, '0' after 8886200 ns,
'1' after 8897000 ns, '0' after 8897050 ns,
'1' after 8907850 ns, '0' after 8907900 ns,
'1' after 8918700 ns, '0' after 8918750 ns,
'1' after 8929550 ns, '0' after 8929600 ns,
'1' after 8940400 ns, '0' after 8940450 ns,
'1' after 8951250 ns, '0' after 8951300 ns,
'1' after 8962100 ns, '0' after 8962150 ns,
'1' after 8972950 ns, '0' after 8973000 ns,
'1' after 8983800 ns, '0' after 8983850 ns,
'1' after 8994650 ns, '0' after 8994700 ns,
'1' after 9005500 ns, '0' after 9005550 ns,
'1' after 9016350 ns, '0' after 9016400 ns,
'1' after 9027200 ns, '0' after 9027250 ns,
'1' after 9038050 ns, '0' after 9038100 ns,
'1' after 9048900 ns, '0' after 9048950 ns,
'1' after 9059750 ns, '0' after 9059800 ns,
'1' after 9070600 ns, '0' after 9070650 ns,
'1' after 9081450 ns, '0' after 9081500 ns,
'1' after 9092300 ns, '0' after 9092350 ns,
'1' after 9103150 ns, '0' after 9103200 ns,
'1' after 9114000 ns, '0' after 9114050 ns,
'1' after 9124850 ns, '0' after 9124900 ns,
'1' after 9135700 ns, '0' after 9135750 ns,
'1' after 9146550 ns, '0' after 9146600 ns,
'1' after 9157400 ns, '0' after 9157450 ns,
'1' after 9168250 ns, '0' after 9168300 ns,
'1' after 9179100 ns, '0' after 9179150 ns,
'1' after 9189950 ns, '0' after 9190000 ns,
'1' after 9200800 ns, '0' after 9200850 ns,
'1' after 9211650 ns, '0' after 9211700 ns,
'1' after 9222500 ns, '0' after 9222550 ns,
'1' after 9233350 ns, '0' after 9233400 ns,
'1' after 9244200 ns, '0' after 9244250 ns,
'1' after 9255050 ns, '0' after 9255100 ns,
'1' after 9265900 ns, '0' after 9265950 ns,
'1' after 9276750 ns, '0' after 9276800 ns,
'1' after 9287600 ns, '0' after 9287650 ns,
'1' after 9298450 ns, '0' after 9298500 ns,
'1' after 9309300 ns, '0' after 9309350 ns,
'1' after 9320150 ns, '0' after 9320200 ns,
'1' after 9331000 ns, '0' after 9331050 ns,
'1' after 9341850 ns, '0' after 9341900 ns,
'1' after 9352700 ns, '0' after 9352750 ns,
'1' after 9363550 ns, '0' after 9363600 ns,
'1' after 9374400 ns, '0' after 9374450 ns,
'1' after 9385250 ns, '0' after 9385300 ns,
'1' after 9396100 ns, '0' after 9396150 ns,
'1' after 9406950 ns, '0' after 9407000 ns,
'1' after 9417800 ns, '0' after 9417850 ns,
'1' after 9428650 ns, '0' after 9428700 ns,
'1' after 9439500 ns, '0' after 9439550 ns,
'1' after 9450350 ns, '0' after 9450400 ns,
'1' after 9461200 ns, '0' after 9461250 ns,
'1' after 9472050 ns, '0' after 9472100 ns,
'1' after 9482900 ns, '0' after 9482950 ns,
'1' after 9493750 ns, '0' after 9493800 ns,
'1' after 9504600 ns, '0' after 9504650 ns,
'1' after 9515450 ns, '0' after 9515500 ns,
'1' after 9526300 ns, '0' after 9526350 ns,
'1' after 9537150 ns, '0' after 9537200 ns,
'1' after 9548000 ns, '0' after 9548050 ns,
'1' after 9558850 ns, '0' after 9558900 ns,
'1' after 9569700 ns, '0' after 9569750 ns,
'1' after 9580550 ns, '0' after 9580600 ns,
'1' after 9591400 ns, '0' after 9591450 ns,
'1' after 9602250 ns, '0' after 9602300 ns,
'1' after 9613100 ns, '0' after 9613150 ns,
'1' after 9623950 ns, '0' after 9624000 ns,
'1' after 9634800 ns, '0' after 9634850 ns,
'1' after 9645650 ns, '0' after 9645700 ns,
'1' after 9656500 ns, '0' after 9656550 ns,
'1' after 9667350 ns, '0' after 9667400 ns,
'1' after 9678200 ns, '0' after 9678250 ns,
'1' after 9689050 ns, '0' after 9689100 ns,
'1' after 9699900 ns, '0' after 9699950 ns,
'1' after 9710750 ns, '0' after 9710800 ns,
'1' after 9721600 ns, '0' after 9721650 ns,
'1' after 9732450 ns, '0' after 9732500 ns,
'1' after 9743300 ns, '0' after 9743350 ns,
'1' after 9754150 ns, '0' after 9754200 ns,
'1' after 9765000 ns, '0' after 9765050 ns,
'1' after 9775850 ns, '0' after 9775900 ns,
'1' after 9786700 ns, '0' after 9786750 ns,
'1' after 9797550 ns, '0' after 9797600 ns,
'1' after 9808400 ns, '0' after 9808450 ns,
'1' after 9819250 ns, '0' after 9819300 ns,
'1' after 9830100 ns, '0' after 9830150 ns,
'1' after 9840950 ns, '0' after 9841000 ns,
'1' after 9851800 ns, '0' after 9851850 ns,
'1' after 9862650 ns, '0' after 9862700 ns,
'1' after 9873500 ns, '0' after 9873550 ns,
'1' after 9884350 ns, '0' after 9884400 ns,
'1' after 9895200 ns, '0' after 9895250 ns,
'1' after 9906050 ns, '0' after 9906100 ns,
'1' after 9916900 ns, '0' after 9916950 ns,
'1' after 9927750 ns, '0' after 9927800 ns,
'1' after 9938600 ns, '0' after 9938650 ns,
'1' after 9949450 ns, '0' after 9949500 ns,
'1' after 9960300 ns, '0' after 9960350 ns,
'1' after 9971150 ns, '0' after 9971200 ns,
'1' after 9982000 ns, '0' after 9982050 ns,
'1' after 9992850 ns, '0' after 9992900 ns,
'1' after 10003700 ns, '0' after 10003750 ns,
'1' after 10014550 ns, '0' after 10014600 ns,
'1' after 10025400 ns, '0' after 10025450 ns,
'1' after 10036250 ns, '0' after 10036300 ns,
'1' after 10047100 ns, '0' after 10047150 ns,
'1' after 10057950 ns, '0' after 10058000 ns,
'1' after 10068800 ns, '0' after 10068850 ns,
'1' after 10079650 ns, '0' after 10079700 ns,
'1' after 10090500 ns, '0' after 10090550 ns,
'1' after 10101350 ns, '0' after 10101400 ns,
'1' after 10112200 ns, '0' after 10112250 ns,
'1' after 10123050 ns, '0' after 10123100 ns,
'1' after 10133900 ns, '0' after 10133950 ns,
'1' after 10144750 ns, '0' after 10144800 ns,
'1' after 10155600 ns, '0' after 10155650 ns,
'1' after 10166450 ns, '0' after 10166500 ns,
'1' after 10177300 ns, '0' after 10177350 ns,
'1' after 10188150 ns, '0' after 10188200 ns,
'1' after 10199000 ns, '0' after 10199050 ns,
'1' after 10209850 ns, '0' after 10209900 ns,
'1' after 10220700 ns, '0' after 10220750 ns,
'1' after 10231550 ns, '0' after 10231600 ns,
'1' after 10242400 ns, '0' after 10242450 ns,
'1' after 10253250 ns, '0' after 10253300 ns,
'1' after 10264100 ns, '0' after 10264150 ns,
'1' after 10274950 ns, '0' after 10275000 ns,
'1' after 10285800 ns, '0' after 10285850 ns,
'1' after 10296650 ns, '0' after 10296700 ns,
'1' after 10307500 ns, '0' after 10307550 ns,
'1' after 10318350 ns, '0' after 10318400 ns,
'1' after 10329200 ns, '0' after 10329250 ns,
'1' after 10340050 ns, '0' after 10340100 ns,
'1' after 10350900 ns, '0' after 10350950 ns,
'1' after 10361750 ns, '0' after 10361800 ns,
'1' after 10372600 ns, '0' after 10372650 ns,
'1' after 10383450 ns, '0' after 10383500 ns,
'1' after 10394300 ns, '0' after 10394350 ns,
'1' after 10405150 ns, '0' after 10405200 ns,
'1' after 10416000 ns, '0' after 10416050 ns,
'1' after 10426850 ns, '0' after 10426900 ns,
'1' after 10437700 ns, '0' after 10437750 ns,
'1' after 10448550 ns, '0' after 10448600 ns,
'1' after 10459400 ns, '0' after 10459450 ns,
'1' after 10470250 ns, '0' after 10470300 ns,
'1' after 10481100 ns, '0' after 10481150 ns,
'1' after 10491950 ns, '0' after 10492000 ns,
'1' after 10502800 ns, '0' after 10502850 ns,
'1' after 10513650 ns, '0' after 10513700 ns,
'1' after 10524500 ns, '0' after 10524550 ns,
'1' after 10535350 ns, '0' after 10535400 ns,
'1' after 10546200 ns, '0' after 10546250 ns,
'1' after 10557050 ns, '0' after 10557100 ns,
'1' after 10567900 ns, '0' after 10567950 ns,
'1' after 10578750 ns, '0' after 10578800 ns,
'1' after 10589600 ns, '0' after 10589650 ns,
'1' after 10600450 ns, '0' after 10600500 ns,
'1' after 10611300 ns, '0' after 10611350 ns,
'1' after 10622150 ns, '0' after 10622200 ns,
'1' after 10633000 ns, '0' after 10633050 ns,
'1' after 10643850 ns, '0' after 10643900 ns,
'1' after 10654700 ns, '0' after 10654750 ns,
'1' after 10665550 ns, '0' after 10665600 ns,
'1' after 10676400 ns, '0' after 10676450 ns,
'1' after 10687250 ns, '0' after 10687300 ns,
'1' after 10698100 ns, '0' after 10698150 ns,
'1' after 10708950 ns, '0' after 10709000 ns,
'1' after 10719800 ns, '0' after 10719850 ns,
'1' after 10730650 ns, '0' after 10730700 ns,
'1' after 10741500 ns, '0' after 10741550 ns,
'1' after 10752350 ns, '0' after 10752400 ns,
'1' after 10763200 ns, '0' after 10763250 ns,
'1' after 10774050 ns, '0' after 10774100 ns,
'1' after 10784900 ns, '0' after 10784950 ns,
'1' after 10795750 ns, '0' after 10795800 ns,
'1' after 10806600 ns, '0' after 10806650 ns,
'1' after 10817450 ns, '0' after 10817500 ns,
'1' after 10828300 ns, '0' after 10828350 ns,
'1' after 10839150 ns, '0' after 10839200 ns,
'1' after 10850000 ns, '0' after 10850050 ns,
'1' after 10860850 ns, '0' after 10860900 ns,
'1' after 10871700 ns, '0' after 10871750 ns,
'1' after 10882550 ns, '0' after 10882600 ns,
'1' after 10893400 ns, '0' after 10893450 ns,
'1' after 10904250 ns, '0' after 10904300 ns,
'1' after 10915100 ns, '0' after 10915150 ns,
'1' after 10925950 ns, '0' after 10926000 ns,
'1' after 10936800 ns, '0' after 10936850 ns,
'1' after 10947650 ns, '0' after 10947700 ns,
'1' after 10958500 ns, '0' after 10958550 ns,
'1' after 10969350 ns, '0' after 10969400 ns,
'1' after 10980200 ns, '0' after 10980250 ns,
'1' after 10991050 ns, '0' after 10991100 ns,
'1' after 11001900 ns, '0' after 11001950 ns,
'1' after 11012750 ns, '0' after 11012800 ns,
'1' after 11023600 ns, '0' after 11023650 ns,
'1' after 11034450 ns, '0' after 11034500 ns,
'1' after 11045300 ns, '0' after 11045350 ns,
'1' after 11056150 ns, '0' after 11056200 ns,
'1' after 11067000 ns, '0' after 11067050 ns,
'1' after 11077850 ns, '0' after 11077900 ns,
'1' after 11088700 ns, '0' after 11088750 ns,
'1' after 11099550 ns, '0' after 11099600 ns,
'1' after 11110400 ns, '0' after 11110450 ns,
'1' after 11121250 ns, '0' after 11121300 ns,
'1' after 11132100 ns, '0' after 11132150 ns,
'1' after 11142950 ns, '0' after 11143000 ns,
'1' after 11153800 ns, '0' after 11153850 ns,
'1' after 11164650 ns, '0' after 11164700 ns,
'1' after 11175500 ns, '0' after 11175550 ns,
'1' after 11186350 ns, '0' after 11186400 ns,
'1' after 11197200 ns, '0' after 11197250 ns,
'1' after 11208050 ns, '0' after 11208100 ns,
'1' after 11218900 ns, '0' after 11218950 ns,
'1' after 11229750 ns, '0' after 11229800 ns,
'1' after 11240600 ns, '0' after 11240650 ns,
'1' after 11251450 ns, '0' after 11251500 ns,
'1' after 11262300 ns, '0' after 11262350 ns,
'1' after 11273150 ns, '0' after 11273200 ns,
'1' after 11284000 ns, '0' after 11284050 ns,
'1' after 11294850 ns, '0' after 11294900 ns,
'1' after 11305700 ns, '0' after 11305750 ns,
'1' after 11316550 ns, '0' after 11316600 ns,
'1' after 11327400 ns, '0' after 11327450 ns,
'1' after 11338250 ns, '0' after 11338300 ns,
'1' after 11349100 ns, '0' after 11349150 ns,
'1' after 11359950 ns, '0' after 11360000 ns,
'1' after 11370800 ns, '0' after 11370850 ns,
'1' after 11381650 ns, '0' after 11381700 ns,
'1' after 11392500 ns, '0' after 11392550 ns,
'1' after 11403350 ns, '0' after 11403400 ns,
'1' after 11414200 ns, '0' after 11414250 ns,
'1' after 11425050 ns, '0' after 11425100 ns,
'1' after 11435900 ns, '0' after 11435950 ns,
'1' after 11446750 ns, '0' after 11446800 ns,
'1' after 11457600 ns, '0' after 11457650 ns,
'1' after 11468450 ns, '0' after 11468500 ns,
'1' after 11479300 ns, '0' after 11479350 ns,
'1' after 11490150 ns, '0' after 11490200 ns,
'1' after 11501000 ns, '0' after 11501050 ns,
'1' after 11511850 ns, '0' after 11511900 ns,
'1' after 11522700 ns, '0' after 11522750 ns,
'1' after 11533550 ns, '0' after 11533600 ns,
'1' after 11544400 ns, '0' after 11544450 ns,
'1' after 11555250 ns, '0' after 11555300 ns,
'1' after 11566100 ns, '0' after 11566150 ns,
'1' after 11576950 ns, '0' after 11577000 ns,
'1' after 11587800 ns, '0' after 11587850 ns,
'1' after 11598650 ns, '0' after 11598700 ns,
'1' after 11609500 ns, '0' after 11609550 ns,
'1' after 11620350 ns, '0' after 11620400 ns,
'1' after 11631200 ns, '0' after 11631250 ns,
'1' after 11642050 ns, '0' after 11642100 ns,
'1' after 11652900 ns, '0' after 11652950 ns,
'1' after 11663750 ns, '0' after 11663800 ns,
'1' after 11674600 ns, '0' after 11674650 ns,
'1' after 11685450 ns, '0' after 11685500 ns,
'1' after 11696300 ns, '0' after 11696350 ns,
'1' after 11707150 ns, '0' after 11707200 ns,
'1' after 11718000 ns, '0' after 11718050 ns,
'1' after 11728850 ns, '0' after 11728900 ns,
'1' after 11739700 ns, '0' after 11739750 ns,
'1' after 11750550 ns, '0' after 11750600 ns,
'1' after 11761400 ns, '0' after 11761450 ns,
'1' after 11772250 ns, '0' after 11772300 ns,
'1' after 11783100 ns, '0' after 11783150 ns,
'1' after 11793950 ns, '0' after 11794000 ns,
'1' after 11804800 ns, '0' after 11804850 ns,
'1' after 11815650 ns, '0' after 11815700 ns,
'1' after 11826500 ns, '0' after 11826550 ns,
'1' after 11837350 ns, '0' after 11837400 ns,
'1' after 11848200 ns, '0' after 11848250 ns,
'1' after 11859050 ns, '0' after 11859100 ns,
'1' after 11869900 ns, '0' after 11869950 ns,
'1' after 11880750 ns, '0' after 11880800 ns,
'1' after 11891600 ns, '0' after 11891650 ns,
'1' after 11902450 ns, '0' after 11902500 ns,
'1' after 11913300 ns, '0' after 11913350 ns,
'1' after 11924150 ns, '0' after 11924200 ns,
'1' after 11935000 ns, '0' after 11935050 ns,
'1' after 11945850 ns, '0' after 11945900 ns,
'1' after 11956700 ns, '0' after 11956750 ns,
'1' after 11967550 ns, '0' after 11967600 ns,
'1' after 11978400 ns, '0' after 11978450 ns,
'1' after 11989250 ns, '0' after 11989300 ns,
'1' after 12000100 ns, '0' after 12000150 ns,
'1' after 12010950 ns, '0' after 12011000 ns,
'1' after 12021800 ns, '0' after 12021850 ns,
'1' after 12032650 ns, '0' after 12032700 ns,
'1' after 12043500 ns, '0' after 12043550 ns,
'1' after 12054350 ns, '0' after 12054400 ns,
'1' after 12065200 ns, '0' after 12065250 ns,
'1' after 12076050 ns, '0' after 12076100 ns,
'1' after 12086900 ns, '0' after 12086950 ns,
'1' after 12097750 ns, '0' after 12097800 ns,
'1' after 12108600 ns, '0' after 12108650 ns,
'1' after 12119450 ns, '0' after 12119500 ns,
'1' after 12130300 ns, '0' after 12130350 ns,
'1' after 12141150 ns, '0' after 12141200 ns,
'1' after 12152000 ns, '0' after 12152050 ns,
'1' after 12162850 ns, '0' after 12162900 ns,
'1' after 12173700 ns, '0' after 12173750 ns,
'1' after 12184550 ns, '0' after 12184600 ns,
'1' after 12195400 ns, '0' after 12195450 ns,
'1' after 12206250 ns, '0' after 12206300 ns,
'1' after 12217100 ns, '0' after 12217150 ns,
'1' after 12227950 ns, '0' after 12228000 ns,
'1' after 12238800 ns, '0' after 12238850 ns,
'1' after 12249650 ns, '0' after 12249700 ns,
'1' after 12260500 ns, '0' after 12260550 ns,
'1' after 12271350 ns, '0' after 12271400 ns,
'1' after 12282200 ns, '0' after 12282250 ns,
'1' after 12293050 ns, '0' after 12293100 ns,
'1' after 12303900 ns, '0' after 12303950 ns,
'1' after 12314750 ns, '0' after 12314800 ns,
'1' after 12325600 ns, '0' after 12325650 ns,
'1' after 12336450 ns, '0' after 12336500 ns,
'1' after 12347300 ns, '0' after 12347350 ns,
'1' after 12358150 ns, '0' after 12358200 ns,
'1' after 12369000 ns, '0' after 12369050 ns,
'1' after 12379850 ns, '0' after 12379900 ns,
'1' after 12390700 ns, '0' after 12390750 ns,
'1' after 12401550 ns, '0' after 12401600 ns,
'1' after 12412400 ns, '0' after 12412450 ns,
'1' after 12423250 ns, '0' after 12423300 ns,
'1' after 12434100 ns, '0' after 12434150 ns,
'1' after 12444950 ns, '0' after 12445000 ns,
'1' after 12455800 ns, '0' after 12455850 ns,
'1' after 12466650 ns, '0' after 12466700 ns,
'1' after 12477500 ns, '0' after 12477550 ns,
'1' after 12488350 ns, '0' after 12488400 ns,
'1' after 12499200 ns, '0' after 12499250 ns,
'1' after 12510050 ns, '0' after 12510100 ns,
'1' after 12520900 ns, '0' after 12520950 ns,
'1' after 12531750 ns, '0' after 12531800 ns,
'1' after 12542600 ns, '0' after 12542650 ns,
'1' after 12553450 ns, '0' after 12553500 ns,
'1' after 12564300 ns, '0' after 12564350 ns,
'1' after 12575150 ns, '0' after 12575200 ns,
'1' after 12586000 ns, '0' after 12586050 ns,
'1' after 12596850 ns, '0' after 12596900 ns,
'1' after 12607700 ns, '0' after 12607750 ns,
'1' after 12618550 ns, '0' after 12618600 ns,
'1' after 12629400 ns, '0' after 12629450 ns,
'1' after 12640250 ns, '0' after 12640300 ns,
'1' after 12651100 ns, '0' after 12651150 ns,
'1' after 12661950 ns, '0' after 12662000 ns,
'1' after 12672800 ns, '0' after 12672850 ns,
'1' after 12683650 ns, '0' after 12683700 ns,
'1' after 12694500 ns, '0' after 12694550 ns,
'1' after 12705350 ns, '0' after 12705400 ns,
'1' after 12716200 ns, '0' after 12716250 ns,
'1' after 12727050 ns, '0' after 12727100 ns,
'1' after 12737900 ns, '0' after 12737950 ns,
'1' after 12748750 ns, '0' after 12748800 ns,
'1' after 12759600 ns, '0' after 12759650 ns,
'1' after 12770450 ns, '0' after 12770500 ns,
'1' after 12781300 ns, '0' after 12781350 ns,
'1' after 12792150 ns, '0' after 12792200 ns,
'1' after 12803000 ns, '0' after 12803050 ns,
'1' after 12813850 ns, '0' after 12813900 ns,
'1' after 12824700 ns, '0' after 12824750 ns,
'1' after 12835550 ns, '0' after 12835600 ns,
'1' after 12846400 ns, '0' after 12846450 ns,
'1' after 12857250 ns, '0' after 12857300 ns,
'1' after 12868100 ns, '0' after 12868150 ns,
'1' after 12878950 ns, '0' after 12879000 ns,
'1' after 12889800 ns, '0' after 12889850 ns,
'1' after 12900650 ns, '0' after 12900700 ns,
'1' after 12911500 ns, '0' after 12911550 ns,
'1' after 12922350 ns, '0' after 12922400 ns,
'1' after 12933200 ns, '0' after 12933250 ns,
'1' after 12944050 ns, '0' after 12944100 ns,
'1' after 12954900 ns, '0' after 12954950 ns,
'1' after 12965750 ns, '0' after 12965800 ns,
'1' after 12976600 ns, '0' after 12976650 ns,
'1' after 12987450 ns, '0' after 12987500 ns,
'1' after 12998300 ns, '0' after 12998350 ns,
'1' after 13009150 ns, '0' after 13009200 ns,
'1' after 13020000 ns, '0' after 13020050 ns,
'1' after 13030850 ns, '0' after 13030900 ns,
'1' after 13041700 ns, '0' after 13041750 ns,
'1' after 13052550 ns, '0' after 13052600 ns,
'1' after 13063400 ns, '0' after 13063450 ns,
'1' after 13074250 ns, '0' after 13074300 ns,
'1' after 13085100 ns, '0' after 13085150 ns,
'1' after 13095950 ns, '0' after 13096000 ns,
'1' after 13106800 ns, '0' after 13106850 ns,
'1' after 13117650 ns, '0' after 13117700 ns,
'1' after 13128500 ns, '0' after 13128550 ns,
'1' after 13139350 ns, '0' after 13139400 ns,
'1' after 13150200 ns, '0' after 13150250 ns,
'1' after 13161050 ns, '0' after 13161100 ns,
'1' after 13171900 ns, '0' after 13171950 ns,
'1' after 13182750 ns, '0' after 13182800 ns,
'1' after 13193600 ns, '0' after 13193650 ns,
'1' after 13204450 ns, '0' after 13204500 ns,
'1' after 13215300 ns, '0' after 13215350 ns,
'1' after 13226150 ns, '0' after 13226200 ns,
'1' after 13237000 ns, '0' after 13237050 ns,
'1' after 13247850 ns, '0' after 13247900 ns,
'1' after 13258700 ns, '0' after 13258750 ns,
'1' after 13269550 ns, '0' after 13269600 ns,
'1' after 13280400 ns, '0' after 13280450 ns,
'1' after 13291250 ns, '0' after 13291300 ns,
'1' after 13302100 ns, '0' after 13302150 ns,
'1' after 13312950 ns, '0' after 13313000 ns,
'1' after 13323800 ns, '0' after 13323850 ns,
'1' after 13334650 ns, '0' after 13334700 ns,
'1' after 13345500 ns, '0' after 13345550 ns,
'1' after 13356350 ns, '0' after 13356400 ns,
'1' after 13367200 ns, '0' after 13367250 ns,
'1' after 13378050 ns, '0' after 13378100 ns,
'1' after 13388900 ns, '0' after 13388950 ns,
'1' after 13399750 ns, '0' after 13399800 ns,
'1' after 13410600 ns, '0' after 13410650 ns,
'1' after 13421450 ns, '0' after 13421500 ns,
'1' after 13432300 ns, '0' after 13432350 ns,
'1' after 13443150 ns, '0' after 13443200 ns,
'1' after 13454000 ns, '0' after 13454050 ns,
'1' after 13464850 ns, '0' after 13464900 ns,
'1' after 13475700 ns, '0' after 13475750 ns,
'1' after 13486550 ns, '0' after 13486600 ns,
'1' after 13497400 ns, '0' after 13497450 ns,
'1' after 13508250 ns, '0' after 13508300 ns,
'1' after 13519100 ns, '0' after 13519150 ns,
'1' after 13529950 ns, '0' after 13530000 ns,
'1' after 13540800 ns, '0' after 13540850 ns,
'1' after 13551650 ns, '0' after 13551700 ns,
'1' after 13562500 ns, '0' after 13562550 ns,
'1' after 13573350 ns, '0' after 13573400 ns,
'1' after 13584200 ns, '0' after 13584250 ns,
'1' after 13595050 ns, '0' after 13595100 ns,
'1' after 13605900 ns, '0' after 13605950 ns,
'1' after 13616750 ns, '0' after 13616800 ns,
'1' after 13627600 ns, '0' after 13627650 ns,
'1' after 13638450 ns, '0' after 13638500 ns,
'1' after 13649300 ns, '0' after 13649350 ns,
'1' after 13660150 ns, '0' after 13660200 ns,
'1' after 13671000 ns, '0' after 13671050 ns,
'1' after 13681850 ns, '0' after 13681900 ns,
'1' after 13692700 ns, '0' after 13692750 ns,
'1' after 13703550 ns, '0' after 13703600 ns,
'1' after 13714400 ns, '0' after 13714450 ns,
'1' after 13725250 ns, '0' after 13725300 ns,
'1' after 13736100 ns, '0' after 13736150 ns,
'1' after 13746950 ns, '0' after 13747000 ns,
'1' after 13757800 ns, '0' after 13757850 ns,
'1' after 13768650 ns, '0' after 13768700 ns,
'1' after 13779500 ns, '0' after 13779550 ns,
'1' after 13790350 ns, '0' after 13790400 ns,
'1' after 13801200 ns, '0' after 13801250 ns,
'1' after 13812050 ns, '0' after 13812100 ns,
'1' after 13822900 ns, '0' after 13822950 ns,
'1' after 13833750 ns, '0' after 13833800 ns,
'1' after 13844600 ns, '0' after 13844650 ns,
'1' after 13855450 ns, '0' after 13855500 ns,
'1' after 13866300 ns, '0' after 13866350 ns,
'1' after 13877150 ns, '0' after 13877200 ns,
'1' after 13888000 ns, '0' after 13888050 ns,
'1' after 13898850 ns, '0' after 13898900 ns,
'1' after 13909700 ns, '0' after 13909750 ns,
'1' after 13920550 ns, '0' after 13920600 ns,
'1' after 13931400 ns, '0' after 13931450 ns,
'1' after 13942250 ns, '0' after 13942300 ns,
'1' after 13953100 ns, '0' after 13953150 ns,
'1' after 13963950 ns, '0' after 13964000 ns,
'1' after 13974800 ns, '0' after 13974850 ns,
'1' after 13985650 ns, '0' after 13985700 ns,
'1' after 13996500 ns, '0' after 13996550 ns,
'1' after 14007350 ns, '0' after 14007400 ns,
'1' after 14018200 ns, '0' after 14018250 ns,
'1' after 14029050 ns, '0' after 14029100 ns,
'1' after 14039900 ns, '0' after 14039950 ns,
'1' after 14050750 ns, '0' after 14050800 ns,
'1' after 14061600 ns, '0' after 14061650 ns,
'1' after 14072450 ns, '0' after 14072500 ns,
'1' after 14083300 ns, '0' after 14083350 ns,
'1' after 14094150 ns, '0' after 14094200 ns,
'1' after 14105000 ns, '0' after 14105050 ns,
'1' after 14115850 ns, '0' after 14115900 ns,
'1' after 14126700 ns, '0' after 14126750 ns,
'1' after 14137550 ns, '0' after 14137600 ns,
'1' after 14148400 ns, '0' after 14148450 ns,
'1' after 14159250 ns, '0' after 14159300 ns,
'1' after 14170100 ns, '0' after 14170150 ns,
'1' after 14180950 ns, '0' after 14181000 ns,
'1' after 14191800 ns, '0' after 14191850 ns,
'1' after 14202650 ns, '0' after 14202700 ns,
'1' after 14213500 ns, '0' after 14213550 ns,
'1' after 14224350 ns, '0' after 14224400 ns,
'1' after 14235200 ns, '0' after 14235250 ns,
'1' after 14246050 ns, '0' after 14246100 ns,
'1' after 14256900 ns, '0' after 14256950 ns,
'1' after 14267750 ns, '0' after 14267800 ns,
'1' after 14278600 ns, '0' after 14278650 ns,
'1' after 14289450 ns, '0' after 14289500 ns,
'1' after 14300300 ns, '0' after 14300350 ns,
'1' after 14311150 ns, '0' after 14311200 ns,
'1' after 14322000 ns, '0' after 14322050 ns,
'1' after 14332850 ns, '0' after 14332900 ns,
'1' after 14343700 ns, '0' after 14343750 ns,
'1' after 14354550 ns, '0' after 14354600 ns,
'1' after 14365400 ns, '0' after 14365450 ns,
'1' after 14376250 ns, '0' after 14376300 ns,
'1' after 14387100 ns, '0' after 14387150 ns,
'1' after 14397950 ns, '0' after 14398000 ns,
'1' after 14408800 ns, '0' after 14408850 ns,
'1' after 14419650 ns, '0' after 14419700 ns,
'1' after 14430500 ns, '0' after 14430550 ns,
'1' after 14441350 ns, '0' after 14441400 ns,
'1' after 14452200 ns, '0' after 14452250 ns,
'1' after 14463050 ns, '0' after 14463100 ns,
'1' after 14473900 ns, '0' after 14473950 ns,
'1' after 14484750 ns, '0' after 14484800 ns,
'1' after 14495600 ns, '0' after 14495650 ns,
'1' after 14506450 ns, '0' after 14506500 ns,
'1' after 14517300 ns, '0' after 14517350 ns,
'1' after 14528150 ns, '0' after 14528200 ns,
'1' after 14539000 ns, '0' after 14539050 ns,
'1' after 14549850 ns, '0' after 14549900 ns,
'1' after 14560700 ns, '0' after 14560750 ns,
'1' after 14571550 ns, '0' after 14571600 ns,
'1' after 14582400 ns, '0' after 14582450 ns,
'1' after 14593250 ns, '0' after 14593300 ns,
'1' after 14604100 ns, '0' after 14604150 ns,
'1' after 14614950 ns, '0' after 14615000 ns,
'1' after 14625800 ns, '0' after 14625850 ns,
'1' after 14636650 ns, '0' after 14636700 ns,
'1' after 14647500 ns, '0' after 14647550 ns,
'1' after 14658350 ns, '0' after 14658400 ns,
'1' after 14669200 ns, '0' after 14669250 ns,
'1' after 14680050 ns, '0' after 14680100 ns,
'1' after 14690900 ns, '0' after 14690950 ns,
'1' after 14701750 ns, '0' after 14701800 ns,
'1' after 14712600 ns, '0' after 14712650 ns,
'1' after 14723450 ns, '0' after 14723500 ns,
'1' after 14734300 ns, '0' after 14734350 ns,
'1' after 14745150 ns, '0' after 14745200 ns,
'1' after 14756000 ns, '0' after 14756050 ns,
'1' after 14766850 ns, '0' after 14766900 ns,
'1' after 14777700 ns, '0' after 14777750 ns,
'1' after 14788550 ns, '0' after 14788600 ns,
'1' after 14799400 ns, '0' after 14799450 ns,
'1' after 14810250 ns, '0' after 14810300 ns,
'1' after 14821100 ns, '0' after 14821150 ns,
'1' after 14831950 ns, '0' after 14832000 ns,
'1' after 14842800 ns, '0' after 14842850 ns,
'1' after 14853650 ns, '0' after 14853700 ns,
'1' after 14864500 ns, '0' after 14864550 ns,
'1' after 14875350 ns, '0' after 14875400 ns,
'1' after 14886200 ns, '0' after 14886250 ns,
'1' after 14897050 ns, '0' after 14897100 ns,
'1' after 14907900 ns, '0' after 14907950 ns,
'1' after 14918750 ns, '0' after 14918800 ns,
'1' after 14929600 ns, '0' after 14929650 ns,
'1' after 14940450 ns, '0' after 14940500 ns,
'1' after 14951300 ns, '0' after 14951350 ns,
'1' after 14962150 ns, '0' after 14962200 ns,
'1' after 14973000 ns, '0' after 14973050 ns,
'1' after 14983850 ns, '0' after 14983900 ns,
'1' after 14994700 ns, '0' after 14994750 ns,
'1' after 15005550 ns, '0' after 15005600 ns,
'1' after 15016400 ns, '0' after 15016450 ns,
'1' after 15027250 ns, '0' after 15027300 ns,
'1' after 15038100 ns, '0' after 15038150 ns,
'1' after 15048950 ns, '0' after 15049000 ns,
'1' after 15059800 ns, '0' after 15059850 ns,
'1' after 15070650 ns, '0' after 15070700 ns,
'1' after 15081500 ns, '0' after 15081550 ns,
'1' after 15092350 ns, '0' after 15092400 ns,
'1' after 15103200 ns, '0' after 15103250 ns,
'1' after 15114050 ns, '0' after 15114100 ns,
'1' after 15124900 ns, '0' after 15124950 ns,
'1' after 15135750 ns, '0' after 15135800 ns,
'1' after 15146600 ns, '0' after 15146650 ns,
'1' after 15157450 ns, '0' after 15157500 ns,
'1' after 15168300 ns, '0' after 15168350 ns,
'1' after 15179150 ns, '0' after 15179200 ns,
'1' after 15190000 ns, '0' after 15190050 ns,
'1' after 15200850 ns, '0' after 15200900 ns,
'1' after 15211700 ns, '0' after 15211750 ns,
'1' after 15222550 ns, '0' after 15222600 ns,
'1' after 15233400 ns, '0' after 15233450 ns,
'1' after 15244250 ns, '0' after 15244300 ns,
'1' after 15255100 ns, '0' after 15255150 ns,
'1' after 15265950 ns, '0' after 15266000 ns,
'1' after 15276800 ns, '0' after 15276850 ns,
'1' after 15287650 ns, '0' after 15287700 ns,
'1' after 15298500 ns, '0' after 15298550 ns,
'1' after 15309350 ns, '0' after 15309400 ns,
'1' after 15320200 ns, '0' after 15320250 ns,
'1' after 15331050 ns, '0' after 15331100 ns,
'1' after 15341900 ns, '0' after 15341950 ns,
'1' after 15352750 ns, '0' after 15352800 ns,
'1' after 15363600 ns, '0' after 15363650 ns,
'1' after 15374450 ns, '0' after 15374500 ns,
'1' after 15385300 ns, '0' after 15385350 ns,
'1' after 15396150 ns, '0' after 15396200 ns,
'1' after 15407000 ns, '0' after 15407050 ns,
'1' after 15417850 ns, '0' after 15417900 ns,
'1' after 15428700 ns, '0' after 15428750 ns,
'1' after 15439550 ns, '0' after 15439600 ns,
'1' after 15450400 ns, '0' after 15450450 ns,
'1' after 15461250 ns, '0' after 15461300 ns,
'1' after 15472100 ns, '0' after 15472150 ns,
'1' after 15482950 ns, '0' after 15483000 ns,
'1' after 15493800 ns, '0' after 15493850 ns,
'1' after 15504650 ns, '0' after 15504700 ns,
'1' after 15515500 ns, '0' after 15515550 ns,
'1' after 15526350 ns, '0' after 15526400 ns,
'1' after 15537200 ns, '0' after 15537250 ns,
'1' after 15548050 ns, '0' after 15548100 ns,
'1' after 15558900 ns, '0' after 15558950 ns,
'1' after 15569750 ns, '0' after 15569800 ns,
'1' after 15580600 ns, '0' after 15580650 ns,
'1' after 15591450 ns, '0' after 15591500 ns,
'1' after 15602300 ns, '0' after 15602350 ns,
'1' after 15613150 ns, '0' after 15613200 ns,
'1' after 15624000 ns, '0' after 15624050 ns,
'1' after 15634850 ns, '0' after 15634900 ns,
'1' after 15645700 ns, '0' after 15645750 ns,
'1' after 15656550 ns, '0' after 15656600 ns,
'1' after 15667400 ns, '0' after 15667450 ns,
'1' after 15678250 ns, '0' after 15678300 ns,
'1' after 15689100 ns, '0' after 15689150 ns,
'1' after 15699950 ns, '0' after 15700000 ns,
'1' after 15710800 ns, '0' after 15710850 ns,
'1' after 15721650 ns, '0' after 15721700 ns,
'1' after 15732500 ns, '0' after 15732550 ns,
'1' after 15743350 ns, '0' after 15743400 ns,
'1' after 15754200 ns, '0' after 15754250 ns,
'1' after 15765050 ns, '0' after 15765100 ns,
'1' after 15775900 ns, '0' after 15775950 ns,
'1' after 15786750 ns, '0' after 15786800 ns,
'1' after 15797600 ns, '0' after 15797650 ns,
'1' after 15808450 ns, '0' after 15808500 ns,
'1' after 15819300 ns, '0' after 15819350 ns,
'1' after 15830150 ns, '0' after 15830200 ns,
'1' after 15841000 ns, '0' after 15841050 ns,
'1' after 15851850 ns, '0' after 15851900 ns,
'1' after 15862700 ns, '0' after 15862750 ns,
'1' after 15873550 ns, '0' after 15873600 ns,
'1' after 15884400 ns, '0' after 15884450 ns,
'1' after 15895250 ns, '0' after 15895300 ns,
'1' after 15906100 ns, '0' after 15906150 ns,
'1' after 15916950 ns, '0' after 15917000 ns,
'1' after 15927800 ns, '0' after 15927850 ns,
'1' after 15938650 ns, '0' after 15938700 ns,
'1' after 15949500 ns, '0' after 15949550 ns,
'1' after 15960350 ns, '0' after 15960400 ns,
'1' after 15971200 ns, '0' after 15971250 ns,
'1' after 15982050 ns, '0' after 15982100 ns,
'1' after 15992900 ns, '0' after 15992950 ns,
'1' after 16003750 ns, '0' after 16003800 ns,
'1' after 16014600 ns, '0' after 16014650 ns,
'1' after 16025450 ns, '0' after 16025500 ns,
'1' after 16036300 ns, '0' after 16036350 ns,
'1' after 16047150 ns, '0' after 16047200 ns,
'1' after 16058000 ns, '0' after 16058050 ns,
'1' after 16068850 ns, '0' after 16068900 ns,
'1' after 16079700 ns, '0' after 16079750 ns,
'1' after 16090550 ns, '0' after 16090600 ns,
'1' after 16101400 ns, '0' after 16101450 ns,
'1' after 16112250 ns, '0' after 16112300 ns,
'1' after 16123100 ns, '0' after 16123150 ns,
'1' after 16133950 ns, '0' after 16134000 ns,
'1' after 16144800 ns, '0' after 16144850 ns,
'1' after 16155650 ns, '0' after 16155700 ns,
'1' after 16166500 ns, '0' after 16166550 ns,
'1' after 16177350 ns, '0' after 16177400 ns,
'1' after 16188200 ns, '0' after 16188250 ns,
'1' after 16199050 ns, '0' after 16199100 ns,
'1' after 16209900 ns, '0' after 16209950 ns,
'1' after 16220750 ns, '0' after 16220800 ns,
'1' after 16231600 ns, '0' after 16231650 ns,
'1' after 16242450 ns, '0' after 16242500 ns,
'1' after 16253300 ns, '0' after 16253350 ns,
'1' after 16264150 ns, '0' after 16264200 ns,
'1' after 16275000 ns, '0' after 16275050 ns,
'1' after 16285850 ns, '0' after 16285900 ns,
'1' after 16296700 ns, '0' after 16296750 ns,
'1' after 16307550 ns, '0' after 16307600 ns,
'1' after 16318400 ns, '0' after 16318450 ns,
'1' after 16329250 ns, '0' after 16329300 ns,
'1' after 16340100 ns, '0' after 16340150 ns,
'1' after 16350950 ns, '0' after 16351000 ns,
'1' after 16361800 ns, '0' after 16361850 ns,
'1' after 16372650 ns, '0' after 16372700 ns,
'1' after 16383500 ns, '0' after 16383550 ns,
'1' after 16394350 ns, '0' after 16394400 ns,
'1' after 16405200 ns, '0' after 16405250 ns,
'1' after 16416050 ns, '0' after 16416100 ns,
'1' after 16426900 ns, '0' after 16426950 ns,
'1' after 16437750 ns, '0' after 16437800 ns,
'1' after 16448600 ns, '0' after 16448650 ns,
'1' after 16459450 ns, '0' after 16459500 ns,
'1' after 16470300 ns, '0' after 16470350 ns,
'1' after 16481150 ns, '0' after 16481200 ns,
'1' after 16492000 ns, '0' after 16492050 ns,
'1' after 16502850 ns, '0' after 16502900 ns,
'1' after 16513700 ns, '0' after 16513750 ns,
'1' after 16524550 ns, '0' after 16524600 ns,
'1' after 16535400 ns, '0' after 16535450 ns,
'1' after 16546250 ns, '0' after 16546300 ns,
'1' after 16557100 ns, '0' after 16557150 ns,
'1' after 16567950 ns, '0' after 16568000 ns,
'1' after 16578800 ns, '0' after 16578850 ns,
'1' after 16589650 ns, '0' after 16589700 ns,
'1' after 16600500 ns, '0' after 16600550 ns,
'1' after 16611350 ns, '0' after 16611400 ns,
'1' after 16622200 ns, '0' after 16622250 ns,
'1' after 16633050 ns, '0' after 16633100 ns,
'1' after 16643900 ns, '0' after 16643950 ns,
'1' after 16654750 ns, '0' after 16654800 ns,
'1' after 16665600 ns, '0' after 16665650 ns,
'1' after 16676450 ns, '0' after 16676500 ns,
'1' after 16687300 ns, '0' after 16687350 ns,
'1' after 16698150 ns, '0' after 16698200 ns,
'1' after 16709000 ns, '0' after 16709050 ns,
'1' after 16719850 ns, '0' after 16719900 ns,
'1' after 16730700 ns, '0' after 16730750 ns,
'1' after 16741550 ns, '0' after 16741600 ns,
'1' after 16752400 ns, '0' after 16752450 ns,
'1' after 16763250 ns, '0' after 16763300 ns,
'1' after 16774100 ns, '0' after 16774150 ns,
'1' after 16784950 ns, '0' after 16785000 ns,
'1' after 16795800 ns, '0' after 16795850 ns,
'1' after 16806650 ns, '0' after 16806700 ns,
'1' after 16817500 ns, '0' after 16817550 ns,
'1' after 16828350 ns, '0' after 16828400 ns,
'1' after 16839200 ns, '0' after 16839250 ns,
'1' after 16850050 ns, '0' after 16850100 ns,
'1' after 16860900 ns, '0' after 16860950 ns,
'1' after 16871750 ns, '0' after 16871800 ns,
'1' after 16882600 ns, '0' after 16882650 ns,
'1' after 16893450 ns, '0' after 16893500 ns,
'1' after 16904300 ns, '0' after 16904350 ns,
'1' after 16915150 ns, '0' after 16915200 ns,
'1' after 16926000 ns, '0' after 16926050 ns,
'1' after 16936850 ns, '0' after 16936900 ns,
'1' after 16947700 ns, '0' after 16947750 ns,
'1' after 16958550 ns, '0' after 16958600 ns,
'1' after 16969400 ns, '0' after 16969450 ns,
'1' after 16980250 ns, '0' after 16980300 ns,
'1' after 16991100 ns, '0' after 16991150 ns,
'1' after 17001950 ns, '0' after 17002000 ns,
'1' after 17012800 ns, '0' after 17012850 ns,
'1' after 17023650 ns, '0' after 17023700 ns,
'1' after 17034500 ns, '0' after 17034550 ns,
'1' after 17045350 ns, '0' after 17045400 ns,
'1' after 17056200 ns, '0' after 17056250 ns,
'1' after 17067050 ns, '0' after 17067100 ns,
'1' after 17077900 ns, '0' after 17077950 ns,
'1' after 17088750 ns, '0' after 17088800 ns,
'1' after 17099600 ns, '0' after 17099650 ns,
'1' after 17110450 ns, '0' after 17110500 ns,
'1' after 17121300 ns, '0' after 17121350 ns,
'1' after 17132150 ns, '0' after 17132200 ns,
'1' after 17143000 ns, '0' after 17143050 ns,
'1' after 17153850 ns, '0' after 17153900 ns,
'1' after 17164700 ns, '0' after 17164750 ns,
'1' after 17175550 ns, '0' after 17175600 ns,
'1' after 17186400 ns, '0' after 17186450 ns,
'1' after 17197250 ns, '0' after 17197300 ns,
'1' after 17208100 ns, '0' after 17208150 ns,
'1' after 17218950 ns, '0' after 17219000 ns,
'1' after 17229800 ns, '0' after 17229850 ns,
'1' after 17240650 ns, '0' after 17240700 ns,
'1' after 17251500 ns, '0' after 17251550 ns,
'1' after 17262350 ns, '0' after 17262400 ns,
'1' after 17273200 ns, '0' after 17273250 ns,
'1' after 17284050 ns, '0' after 17284100 ns,
'1' after 17294900 ns, '0' after 17294950 ns,
'1' after 17305750 ns, '0' after 17305800 ns,
'1' after 17316600 ns, '0' after 17316650 ns,
'1' after 17327450 ns, '0' after 17327500 ns,
'1' after 17338300 ns, '0' after 17338350 ns,
'1' after 17349150 ns, '0' after 17349200 ns,
'1' after 17360000 ns, '0' after 17360050 ns,
'1' after 17370850 ns, '0' after 17370900 ns,
'1' after 17381700 ns, '0' after 17381750 ns,
'1' after 17392550 ns, '0' after 17392600 ns,
'1' after 17403400 ns, '0' after 17403450 ns,
'1' after 17414250 ns, '0' after 17414300 ns,
'1' after 17425100 ns, '0' after 17425150 ns,
'1' after 17435950 ns, '0' after 17436000 ns,
'1' after 17446800 ns, '0' after 17446850 ns,
'1' after 17457650 ns, '0' after 17457700 ns,
'1' after 17468500 ns, '0' after 17468550 ns,
'1' after 17479350 ns, '0' after 17479400 ns,
'1' after 17490200 ns, '0' after 17490250 ns,
'1' after 17501050 ns, '0' after 17501100 ns,
'1' after 17511900 ns, '0' after 17511950 ns,
'1' after 17522750 ns, '0' after 17522800 ns,
'1' after 17533600 ns, '0' after 17533650 ns,
'1' after 17544450 ns, '0' after 17544500 ns,
'1' after 17555300 ns, '0' after 17555350 ns,
'1' after 17566150 ns, '0' after 17566200 ns,
'1' after 17577000 ns, '0' after 17577050 ns,
'1' after 17587850 ns, '0' after 17587900 ns,
'1' after 17598700 ns, '0' after 17598750 ns,
'1' after 17609550 ns, '0' after 17609600 ns,
'1' after 17620400 ns, '0' after 17620450 ns,
'1' after 17631250 ns, '0' after 17631300 ns,
'1' after 17642100 ns, '0' after 17642150 ns,
'1' after 17652950 ns, '0' after 17653000 ns,
'1' after 17663800 ns, '0' after 17663850 ns,
'1' after 17674650 ns, '0' after 17674700 ns,
'1' after 17685500 ns, '0' after 17685550 ns,
'1' after 17696350 ns, '0' after 17696400 ns,
'1' after 17707200 ns, '0' after 17707250 ns,
'1' after 17718050 ns, '0' after 17718100 ns,
'1' after 17728900 ns, '0' after 17728950 ns,
'1' after 17739750 ns, '0' after 17739800 ns,
'1' after 17750600 ns, '0' after 17750650 ns,
'1' after 17761450 ns, '0' after 17761500 ns,
'1' after 17772300 ns, '0' after 17772350 ns,
'1' after 17783150 ns, '0' after 17783200 ns,
'1' after 17794000 ns, '0' after 17794050 ns,
'1' after 17804850 ns, '0' after 17804900 ns,
'1' after 17815700 ns, '0' after 17815750 ns,
'1' after 17826550 ns, '0' after 17826600 ns,
'1' after 17837400 ns, '0' after 17837450 ns,
'1' after 17848250 ns, '0' after 17848300 ns,
'1' after 17859100 ns, '0' after 17859150 ns,
'1' after 17869950 ns, '0' after 17870000 ns,
'1' after 17880800 ns, '0' after 17880850 ns,
'1' after 17891650 ns, '0' after 17891700 ns,
'1' after 17902500 ns, '0' after 17902550 ns,
'1' after 17913350 ns, '0' after 17913400 ns,
'1' after 17924200 ns, '0' after 17924250 ns,
'1' after 17935050 ns, '0' after 17935100 ns,
'1' after 17945900 ns, '0' after 17945950 ns,
'1' after 17956750 ns, '0' after 17956800 ns,
'1' after 17967600 ns, '0' after 17967650 ns,
'1' after 17978450 ns, '0' after 17978500 ns,
'1' after 17989300 ns, '0' after 17989350 ns,
'1' after 18000150 ns, '0' after 18000200 ns,
'1' after 18011000 ns, '0' after 18011050 ns,
'1' after 18021850 ns, '0' after 18021900 ns,
'1' after 18032700 ns, '0' after 18032750 ns,
'1' after 18043550 ns, '0' after 18043600 ns,
'1' after 18054400 ns, '0' after 18054450 ns,
'1' after 18065250 ns, '0' after 18065300 ns,
'1' after 18076100 ns, '0' after 18076150 ns,
'1' after 18086950 ns, '0' after 18087000 ns,
'1' after 18097800 ns, '0' after 18097850 ns,
'1' after 18108650 ns, '0' after 18108700 ns,
'1' after 18119500 ns, '0' after 18119550 ns,
'1' after 18130350 ns, '0' after 18130400 ns,
'1' after 18141200 ns, '0' after 18141250 ns,
'1' after 18152050 ns, '0' after 18152100 ns,
'1' after 18162900 ns, '0' after 18162950 ns,
'1' after 18173750 ns, '0' after 18173800 ns,
'1' after 18184600 ns, '0' after 18184650 ns,
'1' after 18195450 ns, '0' after 18195500 ns,
'1' after 18206300 ns, '0' after 18206350 ns,
'1' after 18217150 ns, '0' after 18217200 ns,
'1' after 18228000 ns, '0' after 18228050 ns,
'1' after 18238850 ns, '0' after 18238900 ns,
'1' after 18249700 ns, '0' after 18249750 ns,
'1' after 18260550 ns, '0' after 18260600 ns,
'1' after 18271400 ns, '0' after 18271450 ns,
'1' after 18282250 ns, '0' after 18282300 ns,
'1' after 18293100 ns, '0' after 18293150 ns,
'1' after 18303950 ns, '0' after 18304000 ns,
'1' after 18314800 ns, '0' after 18314850 ns,
'1' after 18325650 ns, '0' after 18325700 ns,
'1' after 18336500 ns, '0' after 18336550 ns,
'1' after 18347350 ns, '0' after 18347400 ns,
'1' after 18358200 ns, '0' after 18358250 ns,
'1' after 18369050 ns, '0' after 18369100 ns,
'1' after 18379900 ns, '0' after 18379950 ns,
'1' after 18390750 ns, '0' after 18390800 ns,
'1' after 18401600 ns, '0' after 18401650 ns,
'1' after 18412450 ns, '0' after 18412500 ns,
'1' after 18423300 ns, '0' after 18423350 ns,
'1' after 18434150 ns, '0' after 18434200 ns,
'1' after 18445000 ns, '0' after 18445050 ns,
'1' after 18455850 ns, '0' after 18455900 ns,
'1' after 18466700 ns, '0' after 18466750 ns,
'1' after 18477550 ns, '0' after 18477600 ns,
'1' after 18488400 ns, '0' after 18488450 ns,
'1' after 18499250 ns, '0' after 18499300 ns,
'1' after 18510100 ns, '0' after 18510150 ns,
'1' after 18520950 ns, '0' after 18521000 ns,
'1' after 18531800 ns, '0' after 18531850 ns,
'1' after 18542650 ns, '0' after 18542700 ns,
'1' after 18553500 ns, '0' after 18553550 ns,
'1' after 18564350 ns, '0' after 18564400 ns,
'1' after 18575200 ns, '0' after 18575250 ns,
'1' after 18586050 ns, '0' after 18586100 ns,
'1' after 18596900 ns, '0' after 18596950 ns,
'1' after 18607750 ns, '0' after 18607800 ns,
'1' after 18618600 ns, '0' after 18618650 ns,
'1' after 18629450 ns, '0' after 18629500 ns,
'1' after 18640300 ns, '0' after 18640350 ns,
'1' after 18651150 ns, '0' after 18651200 ns,
'1' after 18662000 ns, '0' after 18662050 ns,
'1' after 18672850 ns, '0' after 18672900 ns,
'1' after 18683700 ns, '0' after 18683750 ns,
'1' after 18694550 ns, '0' after 18694600 ns,
'1' after 18705400 ns, '0' after 18705450 ns,
'1' after 18716250 ns, '0' after 18716300 ns,
'1' after 18727100 ns, '0' after 18727150 ns,
'1' after 18737950 ns, '0' after 18738000 ns,
'1' after 18748800 ns, '0' after 18748850 ns,
'1' after 18759650 ns, '0' after 18759700 ns,
'1' after 18770500 ns, '0' after 18770550 ns,
'1' after 18781350 ns, '0' after 18781400 ns,
'1' after 18792200 ns, '0' after 18792250 ns,
'1' after 18803050 ns, '0' after 18803100 ns,
'1' after 18813900 ns, '0' after 18813950 ns,
'1' after 18824750 ns, '0' after 18824800 ns,
'1' after 18835600 ns, '0' after 18835650 ns,
'1' after 18846450 ns, '0' after 18846500 ns,
'1' after 18857300 ns, '0' after 18857350 ns,
'1' after 18868150 ns, '0' after 18868200 ns,
'1' after 18879000 ns, '0' after 18879050 ns,
'1' after 18889850 ns, '0' after 18889900 ns,
'1' after 18900700 ns, '0' after 18900750 ns,
'1' after 18911550 ns, '0' after 18911600 ns,
'1' after 18922400 ns, '0' after 18922450 ns,
'1' after 18933250 ns, '0' after 18933300 ns,
'1' after 18944100 ns, '0' after 18944150 ns,
'1' after 18954950 ns, '0' after 18955000 ns,
'1' after 18965800 ns, '0' after 18965850 ns,
'1' after 18976650 ns, '0' after 18976700 ns,
'1' after 18987500 ns, '0' after 18987550 ns,
'1' after 18998350 ns, '0' after 18998400 ns,
'1' after 19009200 ns, '0' after 19009250 ns,
'1' after 19020050 ns, '0' after 19020100 ns,
'1' after 19030900 ns, '0' after 19030950 ns,
'1' after 19041750 ns, '0' after 19041800 ns,
'1' after 19052600 ns, '0' after 19052650 ns,
'1' after 19063450 ns, '0' after 19063500 ns,
'1' after 19074300 ns, '0' after 19074350 ns,
'1' after 19085150 ns, '0' after 19085200 ns,
'1' after 19096000 ns, '0' after 19096050 ns,
'1' after 19106850 ns, '0' after 19106900 ns,
'1' after 19117700 ns, '0' after 19117750 ns,
'1' after 19128550 ns, '0' after 19128600 ns,
'1' after 19139400 ns, '0' after 19139450 ns,
'1' after 19150250 ns, '0' after 19150300 ns,
'1' after 19161100 ns, '0' after 19161150 ns,
'1' after 19171950 ns, '0' after 19172000 ns,
'1' after 19182800 ns, '0' after 19182850 ns,
'1' after 19193650 ns, '0' after 19193700 ns,
'1' after 19204500 ns, '0' after 19204550 ns,
'1' after 19215350 ns, '0' after 19215400 ns,
'1' after 19226200 ns, '0' after 19226250 ns,
'1' after 19237050 ns, '0' after 19237100 ns,
'1' after 19247900 ns, '0' after 19247950 ns,
'1' after 19258750 ns, '0' after 19258800 ns,
'1' after 19269600 ns, '0' after 19269650 ns,
'1' after 19280450 ns, '0' after 19280500 ns,
'1' after 19291300 ns, '0' after 19291350 ns,
'1' after 19302150 ns, '0' after 19302200 ns,
'1' after 19313000 ns, '0' after 19313050 ns,
'1' after 19323850 ns, '0' after 19323900 ns,
'1' after 19334700 ns, '0' after 19334750 ns,
'1' after 19345550 ns, '0' after 19345600 ns,
'1' after 19356400 ns, '0' after 19356450 ns,
'1' after 19367250 ns, '0' after 19367300 ns,
'1' after 19378100 ns, '0' after 19378150 ns,
'1' after 19388950 ns, '0' after 19389000 ns,
'1' after 19399800 ns, '0' after 19399850 ns,
'1' after 19410650 ns, '0' after 19410700 ns,
'1' after 19421500 ns, '0' after 19421550 ns,
'1' after 19432350 ns, '0' after 19432400 ns,
'1' after 19443200 ns, '0' after 19443250 ns,
'1' after 19454050 ns, '0' after 19454100 ns,
'1' after 19464900 ns, '0' after 19464950 ns,
'1' after 19475750 ns, '0' after 19475800 ns,
'1' after 19486600 ns, '0' after 19486650 ns,
'1' after 19497450 ns, '0' after 19497500 ns,
'1' after 19508300 ns, '0' after 19508350 ns,
'1' after 19519150 ns, '0' after 19519200 ns,
'1' after 19530000 ns, '0' after 19530050 ns,
'1' after 19540850 ns, '0' after 19540900 ns,
'1' after 19551700 ns, '0' after 19551750 ns,
'1' after 19562550 ns, '0' after 19562600 ns,
'1' after 19573400 ns, '0' after 19573450 ns,
'1' after 19584250 ns, '0' after 19584300 ns,
'1' after 19595100 ns, '0' after 19595150 ns,
'1' after 19605950 ns, '0' after 19606000 ns,
'1' after 19616800 ns, '0' after 19616850 ns,
'1' after 19627650 ns, '0' after 19627700 ns,
'1' after 19638500 ns, '0' after 19638550 ns,
'1' after 19649350 ns, '0' after 19649400 ns,
'1' after 19660200 ns, '0' after 19660250 ns,
'1' after 19671050 ns, '0' after 19671100 ns,
'1' after 19681900 ns, '0' after 19681950 ns,
'1' after 19692750 ns, '0' after 19692800 ns,
'1' after 19703600 ns, '0' after 19703650 ns,
'1' after 19714450 ns, '0' after 19714500 ns,
'1' after 19725300 ns, '0' after 19725350 ns,
'1' after 19736150 ns, '0' after 19736200 ns,
'1' after 19747000 ns, '0' after 19747050 ns,
'1' after 19757850 ns, '0' after 19757900 ns,
'1' after 19768700 ns, '0' after 19768750 ns,
'1' after 19779550 ns, '0' after 19779600 ns,
'1' after 19790400 ns, '0' after 19790450 ns,
'1' after 19801250 ns, '0' after 19801300 ns,
'1' after 19812100 ns, '0' after 19812150 ns,
'1' after 19822950 ns, '0' after 19823000 ns,
'1' after 19833800 ns, '0' after 19833850 ns,
'1' after 19844650 ns, '0' after 19844700 ns,
'1' after 19855500 ns, '0' after 19855550 ns,
'1' after 19866350 ns, '0' after 19866400 ns,
'1' after 19877200 ns, '0' after 19877250 ns,
'1' after 19888050 ns, '0' after 19888100 ns,
'1' after 19898900 ns, '0' after 19898950 ns,
'1' after 19909750 ns, '0' after 19909800 ns,
'1' after 19920600 ns, '0' after 19920650 ns,
'1' after 19931450 ns, '0' after 19931500 ns,
'1' after 19942300 ns, '0' after 19942350 ns,
'1' after 19953150 ns, '0' after 19953200 ns,
'1' after 19964000 ns, '0' after 19964050 ns,
'1' after 19974850 ns, '0' after 19974900 ns,
'1' after 19985700 ns, '0' after 19985750 ns,
'1' after 19996550 ns, '0' after 19996600 ns,
'1' after 20007400 ns, '0' after 20007450 ns,
'1' after 20018250 ns, '0' after 20018300 ns,
'1' after 20029100 ns, '0' after 20029150 ns,
'1' after 20039950 ns, '0' after 20040000 ns,
'1' after 20050800 ns, '0' after 20050850 ns,
'1' after 20061650 ns, '0' after 20061700 ns,
'1' after 20072500 ns, '0' after 20072550 ns,
'1' after 20083350 ns, '0' after 20083400 ns,
'1' after 20094200 ns, '0' after 20094250 ns,
'1' after 20105050 ns, '0' after 20105100 ns,
'1' after 20115900 ns, '0' after 20115950 ns,
'1' after 20126750 ns, '0' after 20126800 ns,
'1' after 20137600 ns, '0' after 20137650 ns,
'1' after 20148450 ns, '0' after 20148500 ns,
'1' after 20159300 ns, '0' after 20159350 ns,
'1' after 20170150 ns, '0' after 20170200 ns,
'1' after 20181000 ns, '0' after 20181050 ns,
'1' after 20191850 ns, '0' after 20191900 ns,
'1' after 20202700 ns, '0' after 20202750 ns,
'1' after 20213550 ns, '0' after 20213600 ns,
'1' after 20224400 ns, '0' after 20224450 ns,
'1' after 20235250 ns, '0' after 20235300 ns,
'1' after 20246100 ns, '0' after 20246150 ns,
'1' after 20256950 ns, '0' after 20257000 ns,
'1' after 20267800 ns, '0' after 20267850 ns,
'1' after 20278650 ns, '0' after 20278700 ns,
'1' after 20289500 ns, '0' after 20289550 ns,
'1' after 20300350 ns, '0' after 20300400 ns,
'1' after 20311200 ns, '0' after 20311250 ns,
'1' after 20322050 ns, '0' after 20322100 ns,
'1' after 20332900 ns, '0' after 20332950 ns,
'1' after 20343750 ns, '0' after 20343800 ns,
'1' after 20354600 ns, '0' after 20354650 ns,
'1' after 20365450 ns, '0' after 20365500 ns,
'1' after 20376300 ns, '0' after 20376350 ns,
'1' after 20387150 ns, '0' after 20387200 ns,
'1' after 20398000 ns, '0' after 20398050 ns,
'1' after 20408850 ns, '0' after 20408900 ns,
'1' after 20419700 ns, '0' after 20419750 ns,
'1' after 20430550 ns, '0' after 20430600 ns,
'1' after 20441400 ns, '0' after 20441450 ns,
'1' after 20452250 ns, '0' after 20452300 ns,
'1' after 20463100 ns, '0' after 20463150 ns,
'1' after 20473950 ns, '0' after 20474000 ns,
'1' after 20484800 ns, '0' after 20484850 ns,
'1' after 20495650 ns, '0' after 20495700 ns,
'1' after 20506500 ns, '0' after 20506550 ns,
'1' after 20517350 ns, '0' after 20517400 ns,
'1' after 20528200 ns, '0' after 20528250 ns,
'1' after 20539050 ns, '0' after 20539100 ns,
'1' after 20549900 ns, '0' after 20549950 ns,
'1' after 20560750 ns, '0' after 20560800 ns,
'1' after 20571600 ns, '0' after 20571650 ns,
'1' after 20582450 ns, '0' after 20582500 ns,
'1' after 20593300 ns, '0' after 20593350 ns,
'1' after 20604150 ns, '0' after 20604200 ns,
'1' after 20615000 ns, '0' after 20615050 ns,
'1' after 20625850 ns, '0' after 20625900 ns,
'1' after 20636700 ns, '0' after 20636750 ns,
'1' after 20647550 ns, '0' after 20647600 ns,
'1' after 20658400 ns, '0' after 20658450 ns,
'1' after 20669250 ns, '0' after 20669300 ns,
'1' after 20680100 ns, '0' after 20680150 ns,
'1' after 20690950 ns, '0' after 20691000 ns,
'1' after 20701800 ns, '0' after 20701850 ns,
'1' after 20712650 ns, '0' after 20712700 ns,
'1' after 20723500 ns, '0' after 20723550 ns,
'1' after 20734350 ns, '0' after 20734400 ns,
'1' after 20745200 ns, '0' after 20745250 ns,
'1' after 20756050 ns, '0' after 20756100 ns,
'1' after 20766900 ns, '0' after 20766950 ns,
'1' after 20777750 ns, '0' after 20777800 ns,
'1' after 20788600 ns, '0' after 20788650 ns,
'1' after 20799450 ns, '0' after 20799500 ns,
'1' after 20810300 ns, '0' after 20810350 ns,
'1' after 20821150 ns, '0' after 20821200 ns,
'1' after 20832000 ns, '0' after 20832050 ns,
'1' after 20842850 ns, '0' after 20842900 ns,
'1' after 20853700 ns, '0' after 20853750 ns,
'1' after 20864550 ns, '0' after 20864600 ns,
'1' after 20875400 ns, '0' after 20875450 ns,
'1' after 20886250 ns, '0' after 20886300 ns,
'1' after 20897100 ns, '0' after 20897150 ns,
'1' after 20907950 ns, '0' after 20908000 ns,
'1' after 20918800 ns, '0' after 20918850 ns,
'1' after 20929650 ns, '0' after 20929700 ns,
'1' after 20940500 ns, '0' after 20940550 ns,
'1' after 20951350 ns, '0' after 20951400 ns,
'1' after 20962200 ns, '0' after 20962250 ns,
'1' after 20973050 ns, '0' after 20973100 ns,
'1' after 20983900 ns, '0' after 20983950 ns,
'1' after 20994750 ns, '0' after 20994800 ns,
'1' after 21005600 ns, '0' after 21005650 ns,
'1' after 21016450 ns, '0' after 21016500 ns,
'1' after 21027300 ns, '0' after 21027350 ns,
'1' after 21038150 ns, '0' after 21038200 ns,
'1' after 21049000 ns, '0' after 21049050 ns,
'1' after 21059850 ns, '0' after 21059900 ns,
'1' after 21070700 ns, '0' after 21070750 ns,
'1' after 21081550 ns, '0' after 21081600 ns,
'1' after 21092400 ns, '0' after 21092450 ns,
'1' after 21103250 ns, '0' after 21103300 ns,
'1' after 21114100 ns, '0' after 21114150 ns,
'1' after 21124950 ns, '0' after 21125000 ns,
'1' after 21135800 ns, '0' after 21135850 ns,
'1' after 21146650 ns, '0' after 21146700 ns,
'1' after 21157500 ns, '0' after 21157550 ns,
'1' after 21168350 ns, '0' after 21168400 ns,
'1' after 21179200 ns, '0' after 21179250 ns,
'1' after 21190050 ns, '0' after 21190100 ns,
'1' after 21200900 ns, '0' after 21200950 ns,
'1' after 21211750 ns, '0' after 21211800 ns,
'1' after 21222600 ns, '0' after 21222650 ns,
'1' after 21233450 ns, '0' after 21233500 ns,
'1' after 21244300 ns, '0' after 21244350 ns,
'1' after 21255150 ns, '0' after 21255200 ns,
'1' after 21266000 ns, '0' after 21266050 ns,
'1' after 21276850 ns, '0' after 21276900 ns,
'1' after 21287700 ns, '0' after 21287750 ns,
'1' after 21298550 ns, '0' after 21298600 ns,
'1' after 21309400 ns, '0' after 21309450 ns,
'1' after 21320250 ns, '0' after 21320300 ns,
'1' after 21331100 ns, '0' after 21331150 ns,
'1' after 21341950 ns, '0' after 21342000 ns,
'1' after 21352800 ns, '0' after 21352850 ns,
'1' after 21363650 ns, '0' after 21363700 ns,
'1' after 21374500 ns, '0' after 21374550 ns,
'1' after 21385350 ns, '0' after 21385400 ns,
'1' after 21396200 ns, '0' after 21396250 ns,
'1' after 21407050 ns, '0' after 21407100 ns,
'1' after 21417900 ns, '0' after 21417950 ns,
'1' after 21428750 ns, '0' after 21428800 ns,
'1' after 21439600 ns, '0' after 21439650 ns, -- END OF PROGRAM
'1' after 22201000 ns, '0' after 22201050 ns,
'1' after 22213850 ns, '0' after 22213900 ns, 
'1' after 22224700 ns, '0' after 22224750 ns,
'1' after 22236550 ns, '0' after 22236600 ns;



 -- intr_sig <= '0', '1' after 1000 ns, '0' after 1050 ns;
 -- port_io_sig(30 downto 27) <= "0000", "1000" after 8000 ns;
  --port_io_sig(3 downto 0) <= "1111";
  port_io_sig(30 downto 0) <= (others => 'Z');
  port_io_sig(31) <= '0'; --, '1' after 15000 ns, '0' after 16000 ns;

end architecture behavior;
